// Benchmark "top" written by ABC on Thu May 28 22:01:59 2020

module top ( 
    \in0[0] , \in0[1] , \in0[2] , \in0[3] , \in0[4] , \in0[5] , \in0[6] ,
    \in0[7] , \in0[8] , \in0[9] , \in0[10] , \in0[11] , \in0[12] ,
    \in0[13] , \in0[14] , \in0[15] , \in0[16] , \in0[17] , \in0[18] ,
    \in0[19] , \in0[20] , \in0[21] , \in0[22] , \in0[23] , \in0[24] ,
    \in0[25] , \in0[26] , \in0[27] , \in0[28] , \in0[29] , \in0[30] ,
    \in0[31] , \in0[32] , \in0[33] , \in0[34] , \in0[35] , \in0[36] ,
    \in0[37] , \in0[38] , \in0[39] , \in0[40] , \in0[41] , \in0[42] ,
    \in0[43] , \in0[44] , \in0[45] , \in0[46] , \in0[47] , \in0[48] ,
    \in0[49] , \in0[50] , \in0[51] , \in0[52] , \in0[53] , \in0[54] ,
    \in0[55] , \in0[56] , \in0[57] , \in0[58] , \in0[59] , \in0[60] ,
    \in0[61] , \in0[62] , \in0[63] , \in0[64] , \in0[65] , \in0[66] ,
    \in0[67] , \in0[68] , \in0[69] , \in0[70] , \in0[71] , \in0[72] ,
    \in0[73] , \in0[74] , \in0[75] , \in0[76] , \in0[77] , \in0[78] ,
    \in0[79] , \in0[80] , \in0[81] , \in0[82] , \in0[83] , \in0[84] ,
    \in0[85] , \in0[86] , \in0[87] , \in0[88] , \in0[89] , \in0[90] ,
    \in0[91] , \in0[92] , \in0[93] , \in0[94] , \in0[95] , \in0[96] ,
    \in0[97] , \in0[98] , \in0[99] , \in0[100] , \in0[101] , \in0[102] ,
    \in0[103] , \in0[104] , \in0[105] , \in0[106] , \in0[107] , \in0[108] ,
    \in0[109] , \in0[110] , \in0[111] , \in0[112] , \in0[113] , \in0[114] ,
    \in0[115] , \in0[116] , \in0[117] , \in0[118] , \in0[119] , \in0[120] ,
    \in0[121] , \in0[122] , \in0[123] , \in0[124] , \in0[125] , \in0[126] ,
    \in0[127] , \in1[0] , \in1[1] , \in1[2] , \in1[3] , \in1[4] , \in1[5] ,
    \in1[6] , \in1[7] , \in1[8] , \in1[9] , \in1[10] , \in1[11] ,
    \in1[12] , \in1[13] , \in1[14] , \in1[15] , \in1[16] , \in1[17] ,
    \in1[18] , \in1[19] , \in1[20] , \in1[21] , \in1[22] , \in1[23] ,
    \in1[24] , \in1[25] , \in1[26] , \in1[27] , \in1[28] , \in1[29] ,
    \in1[30] , \in1[31] , \in1[32] , \in1[33] , \in1[34] , \in1[35] ,
    \in1[36] , \in1[37] , \in1[38] , \in1[39] , \in1[40] , \in1[41] ,
    \in1[42] , \in1[43] , \in1[44] , \in1[45] , \in1[46] , \in1[47] ,
    \in1[48] , \in1[49] , \in1[50] , \in1[51] , \in1[52] , \in1[53] ,
    \in1[54] , \in1[55] , \in1[56] , \in1[57] , \in1[58] , \in1[59] ,
    \in1[60] , \in1[61] , \in1[62] , \in1[63] , \in1[64] , \in1[65] ,
    \in1[66] , \in1[67] , \in1[68] , \in1[69] , \in1[70] , \in1[71] ,
    \in1[72] , \in1[73] , \in1[74] , \in1[75] , \in1[76] , \in1[77] ,
    \in1[78] , \in1[79] , \in1[80] , \in1[81] , \in1[82] , \in1[83] ,
    \in1[84] , \in1[85] , \in1[86] , \in1[87] , \in1[88] , \in1[89] ,
    \in1[90] , \in1[91] , \in1[92] , \in1[93] , \in1[94] , \in1[95] ,
    \in1[96] , \in1[97] , \in1[98] , \in1[99] , \in1[100] , \in1[101] ,
    \in1[102] , \in1[103] , \in1[104] , \in1[105] , \in1[106] , \in1[107] ,
    \in1[108] , \in1[109] , \in1[110] , \in1[111] , \in1[112] , \in1[113] ,
    \in1[114] , \in1[115] , \in1[116] , \in1[117] , \in1[118] , \in1[119] ,
    \in1[120] , \in1[121] , \in1[122] , \in1[123] , \in1[124] , \in1[125] ,
    \in1[126] , \in1[127] , \in2[0] , \in2[1] , \in2[2] , \in2[3] ,
    \in2[4] , \in2[5] , \in2[6] , \in2[7] , \in2[8] , \in2[9] , \in2[10] ,
    \in2[11] , \in2[12] , \in2[13] , \in2[14] , \in2[15] , \in2[16] ,
    \in2[17] , \in2[18] , \in2[19] , \in2[20] , \in2[21] , \in2[22] ,
    \in2[23] , \in2[24] , \in2[25] , \in2[26] , \in2[27] , \in2[28] ,
    \in2[29] , \in2[30] , \in2[31] , \in2[32] , \in2[33] , \in2[34] ,
    \in2[35] , \in2[36] , \in2[37] , \in2[38] , \in2[39] , \in2[40] ,
    \in2[41] , \in2[42] , \in2[43] , \in2[44] , \in2[45] , \in2[46] ,
    \in2[47] , \in2[48] , \in2[49] , \in2[50] , \in2[51] , \in2[52] ,
    \in2[53] , \in2[54] , \in2[55] , \in2[56] , \in2[57] , \in2[58] ,
    \in2[59] , \in2[60] , \in2[61] , \in2[62] , \in2[63] , \in2[64] ,
    \in2[65] , \in2[66] , \in2[67] , \in2[68] , \in2[69] , \in2[70] ,
    \in2[71] , \in2[72] , \in2[73] , \in2[74] , \in2[75] , \in2[76] ,
    \in2[77] , \in2[78] , \in2[79] , \in2[80] , \in2[81] , \in2[82] ,
    \in2[83] , \in2[84] , \in2[85] , \in2[86] , \in2[87] , \in2[88] ,
    \in2[89] , \in2[90] , \in2[91] , \in2[92] , \in2[93] , \in2[94] ,
    \in2[95] , \in2[96] , \in2[97] , \in2[98] , \in2[99] , \in2[100] ,
    \in2[101] , \in2[102] , \in2[103] , \in2[104] , \in2[105] , \in2[106] ,
    \in2[107] , \in2[108] , \in2[109] , \in2[110] , \in2[111] , \in2[112] ,
    \in2[113] , \in2[114] , \in2[115] , \in2[116] , \in2[117] , \in2[118] ,
    \in2[119] , \in2[120] , \in2[121] , \in2[122] , \in2[123] , \in2[124] ,
    \in2[125] , \in2[126] , \in2[127] , \in3[0] , \in3[1] , \in3[2] ,
    \in3[3] , \in3[4] , \in3[5] , \in3[6] , \in3[7] , \in3[8] , \in3[9] ,
    \in3[10] , \in3[11] , \in3[12] , \in3[13] , \in3[14] , \in3[15] ,
    \in3[16] , \in3[17] , \in3[18] , \in3[19] , \in3[20] , \in3[21] ,
    \in3[22] , \in3[23] , \in3[24] , \in3[25] , \in3[26] , \in3[27] ,
    \in3[28] , \in3[29] , \in3[30] , \in3[31] , \in3[32] , \in3[33] ,
    \in3[34] , \in3[35] , \in3[36] , \in3[37] , \in3[38] , \in3[39] ,
    \in3[40] , \in3[41] , \in3[42] , \in3[43] , \in3[44] , \in3[45] ,
    \in3[46] , \in3[47] , \in3[48] , \in3[49] , \in3[50] , \in3[51] ,
    \in3[52] , \in3[53] , \in3[54] , \in3[55] , \in3[56] , \in3[57] ,
    \in3[58] , \in3[59] , \in3[60] , \in3[61] , \in3[62] , \in3[63] ,
    \in3[64] , \in3[65] , \in3[66] , \in3[67] , \in3[68] , \in3[69] ,
    \in3[70] , \in3[71] , \in3[72] , \in3[73] , \in3[74] , \in3[75] ,
    \in3[76] , \in3[77] , \in3[78] , \in3[79] , \in3[80] , \in3[81] ,
    \in3[82] , \in3[83] , \in3[84] , \in3[85] , \in3[86] , \in3[87] ,
    \in3[88] , \in3[89] , \in3[90] , \in3[91] , \in3[92] , \in3[93] ,
    \in3[94] , \in3[95] , \in3[96] , \in3[97] , \in3[98] , \in3[99] ,
    \in3[100] , \in3[101] , \in3[102] , \in3[103] , \in3[104] , \in3[105] ,
    \in3[106] , \in3[107] , \in3[108] , \in3[109] , \in3[110] , \in3[111] ,
    \in3[112] , \in3[113] , \in3[114] , \in3[115] , \in3[116] , \in3[117] ,
    \in3[118] , \in3[119] , \in3[120] , \in3[121] , \in3[122] , \in3[123] ,
    \in3[124] , \in3[125] , \in3[126] , \in3[127] ,
    \result[0] , \result[1] , \result[2] , \result[3] , \result[4] ,
    \result[5] , \result[6] , \result[7] , \result[8] , \result[9] ,
    \result[10] , \result[11] , \result[12] , \result[13] , \result[14] ,
    \result[15] , \result[16] , \result[17] , \result[18] , \result[19] ,
    \result[20] , \result[21] , \result[22] , \result[23] , \result[24] ,
    \result[25] , \result[26] , \result[27] , \result[28] , \result[29] ,
    \result[30] , \result[31] , \result[32] , \result[33] , \result[34] ,
    \result[35] , \result[36] , \result[37] , \result[38] , \result[39] ,
    \result[40] , \result[41] , \result[42] , \result[43] , \result[44] ,
    \result[45] , \result[46] , \result[47] , \result[48] , \result[49] ,
    \result[50] , \result[51] , \result[52] , \result[53] , \result[54] ,
    \result[55] , \result[56] , \result[57] , \result[58] , \result[59] ,
    \result[60] , \result[61] , \result[62] , \result[63] , \result[64] ,
    \result[65] , \result[66] , \result[67] , \result[68] , \result[69] ,
    \result[70] , \result[71] , \result[72] , \result[73] , \result[74] ,
    \result[75] , \result[76] , \result[77] , \result[78] , \result[79] ,
    \result[80] , \result[81] , \result[82] , \result[83] , \result[84] ,
    \result[85] , \result[86] , \result[87] , \result[88] , \result[89] ,
    \result[90] , \result[91] , \result[92] , \result[93] , \result[94] ,
    \result[95] , \result[96] , \result[97] , \result[98] , \result[99] ,
    \result[100] , \result[101] , \result[102] , \result[103] ,
    \result[104] , \result[105] , \result[106] , \result[107] ,
    \result[108] , \result[109] , \result[110] , \result[111] ,
    \result[112] , \result[113] , \result[114] , \result[115] ,
    \result[116] , \result[117] , \result[118] , \result[119] ,
    \result[120] , \result[121] , \result[122] , \result[123] ,
    \result[124] , \result[125] , \result[126] , \result[127] ,
    \address[0] , \address[1]   );
  input  \in0[0] , \in0[1] , \in0[2] , \in0[3] , \in0[4] , \in0[5] ,
    \in0[6] , \in0[7] , \in0[8] , \in0[9] , \in0[10] , \in0[11] ,
    \in0[12] , \in0[13] , \in0[14] , \in0[15] , \in0[16] , \in0[17] ,
    \in0[18] , \in0[19] , \in0[20] , \in0[21] , \in0[22] , \in0[23] ,
    \in0[24] , \in0[25] , \in0[26] , \in0[27] , \in0[28] , \in0[29] ,
    \in0[30] , \in0[31] , \in0[32] , \in0[33] , \in0[34] , \in0[35] ,
    \in0[36] , \in0[37] , \in0[38] , \in0[39] , \in0[40] , \in0[41] ,
    \in0[42] , \in0[43] , \in0[44] , \in0[45] , \in0[46] , \in0[47] ,
    \in0[48] , \in0[49] , \in0[50] , \in0[51] , \in0[52] , \in0[53] ,
    \in0[54] , \in0[55] , \in0[56] , \in0[57] , \in0[58] , \in0[59] ,
    \in0[60] , \in0[61] , \in0[62] , \in0[63] , \in0[64] , \in0[65] ,
    \in0[66] , \in0[67] , \in0[68] , \in0[69] , \in0[70] , \in0[71] ,
    \in0[72] , \in0[73] , \in0[74] , \in0[75] , \in0[76] , \in0[77] ,
    \in0[78] , \in0[79] , \in0[80] , \in0[81] , \in0[82] , \in0[83] ,
    \in0[84] , \in0[85] , \in0[86] , \in0[87] , \in0[88] , \in0[89] ,
    \in0[90] , \in0[91] , \in0[92] , \in0[93] , \in0[94] , \in0[95] ,
    \in0[96] , \in0[97] , \in0[98] , \in0[99] , \in0[100] , \in0[101] ,
    \in0[102] , \in0[103] , \in0[104] , \in0[105] , \in0[106] , \in0[107] ,
    \in0[108] , \in0[109] , \in0[110] , \in0[111] , \in0[112] , \in0[113] ,
    \in0[114] , \in0[115] , \in0[116] , \in0[117] , \in0[118] , \in0[119] ,
    \in0[120] , \in0[121] , \in0[122] , \in0[123] , \in0[124] , \in0[125] ,
    \in0[126] , \in0[127] , \in1[0] , \in1[1] , \in1[2] , \in1[3] ,
    \in1[4] , \in1[5] , \in1[6] , \in1[7] , \in1[8] , \in1[9] , \in1[10] ,
    \in1[11] , \in1[12] , \in1[13] , \in1[14] , \in1[15] , \in1[16] ,
    \in1[17] , \in1[18] , \in1[19] , \in1[20] , \in1[21] , \in1[22] ,
    \in1[23] , \in1[24] , \in1[25] , \in1[26] , \in1[27] , \in1[28] ,
    \in1[29] , \in1[30] , \in1[31] , \in1[32] , \in1[33] , \in1[34] ,
    \in1[35] , \in1[36] , \in1[37] , \in1[38] , \in1[39] , \in1[40] ,
    \in1[41] , \in1[42] , \in1[43] , \in1[44] , \in1[45] , \in1[46] ,
    \in1[47] , \in1[48] , \in1[49] , \in1[50] , \in1[51] , \in1[52] ,
    \in1[53] , \in1[54] , \in1[55] , \in1[56] , \in1[57] , \in1[58] ,
    \in1[59] , \in1[60] , \in1[61] , \in1[62] , \in1[63] , \in1[64] ,
    \in1[65] , \in1[66] , \in1[67] , \in1[68] , \in1[69] , \in1[70] ,
    \in1[71] , \in1[72] , \in1[73] , \in1[74] , \in1[75] , \in1[76] ,
    \in1[77] , \in1[78] , \in1[79] , \in1[80] , \in1[81] , \in1[82] ,
    \in1[83] , \in1[84] , \in1[85] , \in1[86] , \in1[87] , \in1[88] ,
    \in1[89] , \in1[90] , \in1[91] , \in1[92] , \in1[93] , \in1[94] ,
    \in1[95] , \in1[96] , \in1[97] , \in1[98] , \in1[99] , \in1[100] ,
    \in1[101] , \in1[102] , \in1[103] , \in1[104] , \in1[105] , \in1[106] ,
    \in1[107] , \in1[108] , \in1[109] , \in1[110] , \in1[111] , \in1[112] ,
    \in1[113] , \in1[114] , \in1[115] , \in1[116] , \in1[117] , \in1[118] ,
    \in1[119] , \in1[120] , \in1[121] , \in1[122] , \in1[123] , \in1[124] ,
    \in1[125] , \in1[126] , \in1[127] , \in2[0] , \in2[1] , \in2[2] ,
    \in2[3] , \in2[4] , \in2[5] , \in2[6] , \in2[7] , \in2[8] , \in2[9] ,
    \in2[10] , \in2[11] , \in2[12] , \in2[13] , \in2[14] , \in2[15] ,
    \in2[16] , \in2[17] , \in2[18] , \in2[19] , \in2[20] , \in2[21] ,
    \in2[22] , \in2[23] , \in2[24] , \in2[25] , \in2[26] , \in2[27] ,
    \in2[28] , \in2[29] , \in2[30] , \in2[31] , \in2[32] , \in2[33] ,
    \in2[34] , \in2[35] , \in2[36] , \in2[37] , \in2[38] , \in2[39] ,
    \in2[40] , \in2[41] , \in2[42] , \in2[43] , \in2[44] , \in2[45] ,
    \in2[46] , \in2[47] , \in2[48] , \in2[49] , \in2[50] , \in2[51] ,
    \in2[52] , \in2[53] , \in2[54] , \in2[55] , \in2[56] , \in2[57] ,
    \in2[58] , \in2[59] , \in2[60] , \in2[61] , \in2[62] , \in2[63] ,
    \in2[64] , \in2[65] , \in2[66] , \in2[67] , \in2[68] , \in2[69] ,
    \in2[70] , \in2[71] , \in2[72] , \in2[73] , \in2[74] , \in2[75] ,
    \in2[76] , \in2[77] , \in2[78] , \in2[79] , \in2[80] , \in2[81] ,
    \in2[82] , \in2[83] , \in2[84] , \in2[85] , \in2[86] , \in2[87] ,
    \in2[88] , \in2[89] , \in2[90] , \in2[91] , \in2[92] , \in2[93] ,
    \in2[94] , \in2[95] , \in2[96] , \in2[97] , \in2[98] , \in2[99] ,
    \in2[100] , \in2[101] , \in2[102] , \in2[103] , \in2[104] , \in2[105] ,
    \in2[106] , \in2[107] , \in2[108] , \in2[109] , \in2[110] , \in2[111] ,
    \in2[112] , \in2[113] , \in2[114] , \in2[115] , \in2[116] , \in2[117] ,
    \in2[118] , \in2[119] , \in2[120] , \in2[121] , \in2[122] , \in2[123] ,
    \in2[124] , \in2[125] , \in2[126] , \in2[127] , \in3[0] , \in3[1] ,
    \in3[2] , \in3[3] , \in3[4] , \in3[5] , \in3[6] , \in3[7] , \in3[8] ,
    \in3[9] , \in3[10] , \in3[11] , \in3[12] , \in3[13] , \in3[14] ,
    \in3[15] , \in3[16] , \in3[17] , \in3[18] , \in3[19] , \in3[20] ,
    \in3[21] , \in3[22] , \in3[23] , \in3[24] , \in3[25] , \in3[26] ,
    \in3[27] , \in3[28] , \in3[29] , \in3[30] , \in3[31] , \in3[32] ,
    \in3[33] , \in3[34] , \in3[35] , \in3[36] , \in3[37] , \in3[38] ,
    \in3[39] , \in3[40] , \in3[41] , \in3[42] , \in3[43] , \in3[44] ,
    \in3[45] , \in3[46] , \in3[47] , \in3[48] , \in3[49] , \in3[50] ,
    \in3[51] , \in3[52] , \in3[53] , \in3[54] , \in3[55] , \in3[56] ,
    \in3[57] , \in3[58] , \in3[59] , \in3[60] , \in3[61] , \in3[62] ,
    \in3[63] , \in3[64] , \in3[65] , \in3[66] , \in3[67] , \in3[68] ,
    \in3[69] , \in3[70] , \in3[71] , \in3[72] , \in3[73] , \in3[74] ,
    \in3[75] , \in3[76] , \in3[77] , \in3[78] , \in3[79] , \in3[80] ,
    \in3[81] , \in3[82] , \in3[83] , \in3[84] , \in3[85] , \in3[86] ,
    \in3[87] , \in3[88] , \in3[89] , \in3[90] , \in3[91] , \in3[92] ,
    \in3[93] , \in3[94] , \in3[95] , \in3[96] , \in3[97] , \in3[98] ,
    \in3[99] , \in3[100] , \in3[101] , \in3[102] , \in3[103] , \in3[104] ,
    \in3[105] , \in3[106] , \in3[107] , \in3[108] , \in3[109] , \in3[110] ,
    \in3[111] , \in3[112] , \in3[113] , \in3[114] , \in3[115] , \in3[116] ,
    \in3[117] , \in3[118] , \in3[119] , \in3[120] , \in3[121] , \in3[122] ,
    \in3[123] , \in3[124] , \in3[125] , \in3[126] , \in3[127] ;
  output \result[0] , \result[1] , \result[2] , \result[3] , \result[4] ,
    \result[5] , \result[6] , \result[7] , \result[8] , \result[9] ,
    \result[10] , \result[11] , \result[12] , \result[13] , \result[14] ,
    \result[15] , \result[16] , \result[17] , \result[18] , \result[19] ,
    \result[20] , \result[21] , \result[22] , \result[23] , \result[24] ,
    \result[25] , \result[26] , \result[27] , \result[28] , \result[29] ,
    \result[30] , \result[31] , \result[32] , \result[33] , \result[34] ,
    \result[35] , \result[36] , \result[37] , \result[38] , \result[39] ,
    \result[40] , \result[41] , \result[42] , \result[43] , \result[44] ,
    \result[45] , \result[46] , \result[47] , \result[48] , \result[49] ,
    \result[50] , \result[51] , \result[52] , \result[53] , \result[54] ,
    \result[55] , \result[56] , \result[57] , \result[58] , \result[59] ,
    \result[60] , \result[61] , \result[62] , \result[63] , \result[64] ,
    \result[65] , \result[66] , \result[67] , \result[68] , \result[69] ,
    \result[70] , \result[71] , \result[72] , \result[73] , \result[74] ,
    \result[75] , \result[76] , \result[77] , \result[78] , \result[79] ,
    \result[80] , \result[81] , \result[82] , \result[83] , \result[84] ,
    \result[85] , \result[86] , \result[87] , \result[88] , \result[89] ,
    \result[90] , \result[91] , \result[92] , \result[93] , \result[94] ,
    \result[95] , \result[96] , \result[97] , \result[98] , \result[99] ,
    \result[100] , \result[101] , \result[102] , \result[103] ,
    \result[104] , \result[105] , \result[106] , \result[107] ,
    \result[108] , \result[109] , \result[110] , \result[111] ,
    \result[112] , \result[113] , \result[114] , \result[115] ,
    \result[116] , \result[117] , \result[118] , \result[119] ,
    \result[120] , \result[121] , \result[122] , \result[123] ,
    \result[124] , \result[125] , \result[126] , \result[127] ,
    \address[0] , \address[1] ;
  wire n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
    n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
    n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
    n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
    n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
    n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
    n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
    n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
    n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
    n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
    n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
    n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
    n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
    n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
    n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
    n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
    n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
    n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
    n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
    n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
    n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
    n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
    n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
    n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
    n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
    n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
    n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
    n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
    n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
    n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
    n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
    n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
    n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
    n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
    n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
    n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
    n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
    n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
    n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
    n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
    n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
    n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
    n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
    n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
    n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
    n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
    n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
    n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
    n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
    n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
    n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
    n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
    n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
    n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
    n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
    n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
    n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
    n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
    n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
    n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
    n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
    n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
    n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
    n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
    n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
    n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
    n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
    n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
    n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
    n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
    n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409,
    n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419,
    n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429,
    n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439,
    n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449,
    n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459,
    n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469,
    n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479,
    n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489,
    n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499,
    n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509,
    n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519,
    n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529,
    n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539,
    n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549,
    n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559,
    n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569,
    n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579,
    n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589,
    n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599,
    n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609,
    n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619,
    n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629,
    n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639,
    n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649,
    n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659,
    n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669,
    n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679,
    n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689,
    n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699,
    n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709,
    n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719,
    n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729,
    n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739,
    n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749,
    n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759,
    n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769,
    n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779,
    n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789,
    n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799,
    n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809,
    n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819,
    n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829,
    n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839,
    n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849,
    n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859,
    n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869,
    n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879,
    n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889,
    n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899,
    n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909,
    n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919,
    n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929,
    n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939,
    n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949,
    n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959,
    n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969,
    n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979,
    n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989,
    n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999,
    n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009,
    n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019,
    n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029,
    n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039,
    n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049,
    n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059,
    n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069,
    n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079,
    n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089,
    n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099,
    n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109,
    n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119,
    n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129,
    n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139,
    n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149,
    n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159,
    n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169,
    n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179,
    n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189,
    n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199,
    n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209,
    n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219,
    n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229,
    n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239,
    n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249,
    n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259,
    n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269,
    n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279,
    n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289,
    n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299,
    n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309,
    n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319,
    n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329,
    n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339,
    n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349,
    n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359,
    n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369,
    n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379,
    n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389,
    n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399,
    n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409,
    n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419,
    n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429,
    n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439,
    n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449,
    n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459,
    n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469,
    n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479,
    n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489,
    n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499,
    n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509,
    n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519,
    n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529,
    n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539,
    n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549,
    n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559,
    n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569,
    n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579,
    n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589,
    n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599,
    n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609,
    n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619,
    n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629,
    n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639,
    n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649,
    n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659,
    n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669,
    n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679,
    n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689,
    n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699,
    n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709,
    n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719,
    n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729,
    n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739,
    n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749,
    n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759,
    n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769,
    n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779,
    n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789,
    n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799,
    n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809,
    n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819,
    n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829,
    n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839,
    n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849,
    n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859,
    n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869,
    n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879,
    n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889,
    n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899,
    n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909,
    n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919,
    n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929,
    n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939,
    n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949,
    n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959,
    n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969,
    n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979,
    n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989,
    n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999,
    n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009,
    n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019,
    n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029,
    n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039,
    n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049,
    n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059,
    n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069,
    n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079,
    n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089,
    n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099,
    n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109,
    n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119,
    n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129,
    n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139,
    n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149,
    n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159,
    n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169,
    n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179,
    n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189,
    n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199,
    n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209,
    n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219,
    n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229,
    n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239,
    n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249,
    n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259,
    n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269,
    n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279,
    n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289,
    n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299,
    n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309,
    n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319,
    n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329,
    n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339,
    n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349,
    n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359,
    n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369,
    n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379,
    n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389,
    n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399,
    n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409,
    n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419,
    n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429,
    n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439,
    n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449,
    n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459,
    n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469,
    n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479,
    n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489,
    n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499,
    n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509,
    n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519,
    n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529,
    n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539,
    n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549,
    n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559,
    n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569,
    n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579,
    n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589,
    n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599,
    n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609,
    n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619,
    n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629,
    n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639,
    n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649,
    n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659,
    n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669,
    n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679,
    n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689,
    n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699,
    n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709,
    n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719,
    n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729,
    n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739,
    n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749,
    n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759,
    n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769,
    n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779,
    n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789,
    n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799,
    n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809,
    n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819,
    n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829,
    n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839,
    n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849,
    n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859,
    n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869,
    n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879,
    n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889,
    n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899,
    n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909,
    n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919,
    n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929,
    n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939,
    n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949,
    n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959,
    n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969,
    n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979,
    n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989,
    n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999,
    n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009,
    n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019,
    n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029,
    n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039,
    n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049,
    n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059,
    n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069,
    n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079,
    n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089,
    n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099,
    n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109,
    n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119,
    n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129,
    n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139,
    n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149,
    n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159,
    n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169,
    n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179,
    n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189,
    n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199,
    n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209,
    n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219,
    n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229,
    n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239,
    n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249,
    n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259,
    n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269,
    n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280,
    n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290,
    n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300,
    n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310,
    n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320,
    n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330,
    n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340,
    n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350,
    n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360,
    n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370,
    n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380,
    n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390,
    n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400,
    n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410,
    n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420,
    n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430,
    n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440,
    n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450,
    n4451, n4452, n4453, n4455, n4456, n4458, n4459, n4461, n4462, n4464,
    n4465, n4467, n4468, n4470, n4471, n4473, n4474, n4476, n4477, n4479,
    n4480, n4482, n4483, n4485, n4486, n4488, n4489, n4491, n4492, n4494,
    n4495, n4497, n4498, n4500, n4501, n4503, n4504, n4506, n4507, n4509,
    n4510, n4512, n4513, n4515, n4516, n4518, n4519, n4521, n4522, n4524,
    n4525, n4527, n4528, n4530, n4531, n4533, n4534, n4536, n4537, n4539,
    n4540, n4542, n4543, n4545, n4546, n4548, n4549, n4551, n4552, n4554,
    n4555, n4557, n4558, n4560, n4561, n4563, n4564, n4566, n4567, n4569,
    n4570, n4572, n4573, n4575, n4576, n4578, n4579, n4581, n4582, n4584,
    n4585, n4587, n4588, n4590, n4591, n4593, n4594, n4596, n4597, n4599,
    n4600, n4602, n4603, n4605, n4606, n4608, n4609, n4611, n4612, n4614,
    n4615, n4617, n4618, n4620, n4621, n4623, n4624, n4626, n4627, n4629,
    n4630, n4632, n4633, n4635, n4636, n4638, n4639, n4641, n4642, n4644,
    n4645, n4647, n4648, n4650, n4651, n4653, n4654, n4656, n4657, n4659,
    n4660, n4662, n4663, n4665, n4666, n4668, n4669, n4671, n4672, n4674,
    n4675, n4677, n4678, n4680, n4681, n4683, n4684, n4686, n4687, n4689,
    n4690, n4692, n4693, n4695, n4696, n4698, n4699, n4701, n4702, n4704,
    n4705, n4707, n4708, n4710, n4711, n4713, n4714, n4716, n4717, n4719,
    n4720, n4722, n4723, n4725, n4726, n4728, n4729, n4731, n4732, n4734,
    n4735, n4737, n4738, n4740, n4741, n4743, n4744, n4746, n4747, n4749,
    n4750, n4752, n4753, n4755, n4756, n4758, n4759, n4761, n4762, n4764,
    n4765, n4767, n4768, n4770, n4771, n4773, n4774, n4776, n4777, n4779,
    n4780, n4782, n4783, n4785, n4786, n4788, n4789, n4791, n4792, n4794,
    n4795, n4797, n4798, n4800, n4801, n4803, n4804, n4806, n4807, n4809,
    n4810, n4812, n4813, n4815, n4816, n4818, n4819, n4821, n4822, n4824,
    n4825, n4827, n4828, n4830, n4831, n4834, n4835;
  jnot g0000(.din(\in2[30] ), .dout(n642));
  jand g0001(.dina(\in3[30] ), .dinb(n642), .dout(n643));
  jnot g0002(.din(n643), .dout(n644));
  jnot g0003(.din(\in3[29] ), .dout(n645));
  jand g0004(.dina(n645), .dinb(\in2[29] ), .dout(n646));
  jnot g0005(.din(\in2[29] ), .dout(n647));
  jand g0006(.dina(\in3[29] ), .dinb(n647), .dout(n648));
  jnot g0007(.din(n648), .dout(n649));
  jnot g0008(.din(\in3[28] ), .dout(n650));
  jand g0009(.dina(n650), .dinb(\in2[28] ), .dout(n651));
  jnot g0010(.din(\in2[28] ), .dout(n652));
  jand g0011(.dina(\in3[28] ), .dinb(n652), .dout(n653));
  jnot g0012(.din(n653), .dout(n654));
  jnot g0013(.din(\in3[27] ), .dout(n655));
  jand g0014(.dina(n655), .dinb(\in2[27] ), .dout(n656));
  jnot g0015(.din(\in2[27] ), .dout(n657));
  jand g0016(.dina(\in3[27] ), .dinb(n657), .dout(n658));
  jnot g0017(.din(n658), .dout(n659));
  jnot g0018(.din(\in3[26] ), .dout(n660));
  jand g0019(.dina(n660), .dinb(\in2[26] ), .dout(n661));
  jnot g0020(.din(\in2[26] ), .dout(n662));
  jand g0021(.dina(\in3[26] ), .dinb(n662), .dout(n663));
  jnot g0022(.din(n663), .dout(n664));
  jnot g0023(.din(\in3[25] ), .dout(n665));
  jand g0024(.dina(n665), .dinb(\in2[25] ), .dout(n666));
  jnot g0025(.din(\in2[25] ), .dout(n667));
  jand g0026(.dina(\in3[25] ), .dinb(n667), .dout(n668));
  jnot g0027(.din(n668), .dout(n669));
  jnot g0028(.din(\in3[24] ), .dout(n670));
  jand g0029(.dina(n670), .dinb(\in2[24] ), .dout(n671));
  jnot g0030(.din(\in2[24] ), .dout(n672));
  jand g0031(.dina(\in3[24] ), .dinb(n672), .dout(n673));
  jnot g0032(.din(n673), .dout(n674));
  jnot g0033(.din(\in3[23] ), .dout(n675));
  jand g0034(.dina(n675), .dinb(\in2[23] ), .dout(n676));
  jnot g0035(.din(\in2[23] ), .dout(n677));
  jand g0036(.dina(\in3[23] ), .dinb(n677), .dout(n678));
  jnot g0037(.din(n678), .dout(n679));
  jnot g0038(.din(\in3[22] ), .dout(n680));
  jand g0039(.dina(n680), .dinb(\in2[22] ), .dout(n681));
  jnot g0040(.din(\in2[22] ), .dout(n682));
  jand g0041(.dina(\in3[22] ), .dinb(n682), .dout(n683));
  jnot g0042(.din(n683), .dout(n684));
  jnot g0043(.din(\in3[21] ), .dout(n685));
  jand g0044(.dina(n685), .dinb(\in2[21] ), .dout(n686));
  jnot g0045(.din(\in2[21] ), .dout(n687));
  jand g0046(.dina(\in3[21] ), .dinb(n687), .dout(n688));
  jnot g0047(.din(n688), .dout(n689));
  jnot g0048(.din(\in3[20] ), .dout(n690));
  jand g0049(.dina(n690), .dinb(\in2[20] ), .dout(n691));
  jnot g0050(.din(\in2[20] ), .dout(n692));
  jand g0051(.dina(\in3[20] ), .dinb(n692), .dout(n693));
  jnot g0052(.din(n693), .dout(n694));
  jnot g0053(.din(\in3[19] ), .dout(n695));
  jand g0054(.dina(n695), .dinb(\in2[19] ), .dout(n696));
  jnot g0055(.din(\in2[19] ), .dout(n697));
  jand g0056(.dina(\in3[19] ), .dinb(n697), .dout(n698));
  jnot g0057(.din(n698), .dout(n699));
  jnot g0058(.din(\in3[18] ), .dout(n700));
  jand g0059(.dina(n700), .dinb(\in2[18] ), .dout(n701));
  jnot g0060(.din(\in2[18] ), .dout(n702));
  jand g0061(.dina(\in3[18] ), .dinb(n702), .dout(n703));
  jnot g0062(.din(n703), .dout(n704));
  jnot g0063(.din(\in3[17] ), .dout(n705));
  jand g0064(.dina(n705), .dinb(\in2[17] ), .dout(n706));
  jnot g0065(.din(\in2[17] ), .dout(n707));
  jand g0066(.dina(\in3[17] ), .dinb(n707), .dout(n708));
  jnot g0067(.din(n708), .dout(n709));
  jnot g0068(.din(\in3[16] ), .dout(n710));
  jand g0069(.dina(n710), .dinb(\in2[16] ), .dout(n711));
  jnot g0070(.din(\in2[16] ), .dout(n712));
  jand g0071(.dina(\in3[16] ), .dinb(n712), .dout(n713));
  jnot g0072(.din(n713), .dout(n714));
  jnot g0073(.din(\in3[15] ), .dout(n715));
  jand g0074(.dina(n715), .dinb(\in2[15] ), .dout(n716));
  jnot g0075(.din(\in2[15] ), .dout(n717));
  jand g0076(.dina(\in3[15] ), .dinb(n717), .dout(n718));
  jnot g0077(.din(n718), .dout(n719));
  jnot g0078(.din(\in3[14] ), .dout(n720));
  jand g0079(.dina(n720), .dinb(\in2[14] ), .dout(n721));
  jnot g0080(.din(\in2[14] ), .dout(n722));
  jand g0081(.dina(\in3[14] ), .dinb(n722), .dout(n723));
  jnot g0082(.din(n723), .dout(n724));
  jnot g0083(.din(\in3[13] ), .dout(n725));
  jand g0084(.dina(n725), .dinb(\in2[13] ), .dout(n726));
  jnot g0085(.din(\in2[13] ), .dout(n727));
  jand g0086(.dina(\in3[13] ), .dinb(n727), .dout(n728));
  jnot g0087(.din(n728), .dout(n729));
  jnot g0088(.din(\in3[12] ), .dout(n730));
  jand g0089(.dina(n730), .dinb(\in2[12] ), .dout(n731));
  jnot g0090(.din(\in2[12] ), .dout(n732));
  jand g0091(.dina(\in3[12] ), .dinb(n732), .dout(n733));
  jnot g0092(.din(n733), .dout(n734));
  jnot g0093(.din(\in3[11] ), .dout(n735));
  jand g0094(.dina(n735), .dinb(\in2[11] ), .dout(n736));
  jnot g0095(.din(\in2[11] ), .dout(n737));
  jand g0096(.dina(\in3[11] ), .dinb(n737), .dout(n738));
  jnot g0097(.din(n738), .dout(n739));
  jnot g0098(.din(\in3[10] ), .dout(n740));
  jand g0099(.dina(n740), .dinb(\in2[10] ), .dout(n741));
  jnot g0100(.din(\in2[10] ), .dout(n742));
  jand g0101(.dina(\in3[10] ), .dinb(n742), .dout(n743));
  jnot g0102(.din(n743), .dout(n744));
  jnot g0103(.din(\in3[9] ), .dout(n745));
  jand g0104(.dina(n745), .dinb(\in2[9] ), .dout(n746));
  jnot g0105(.din(\in2[9] ), .dout(n747));
  jand g0106(.dina(\in3[9] ), .dinb(n747), .dout(n748));
  jnot g0107(.din(n748), .dout(n749));
  jnot g0108(.din(\in3[8] ), .dout(n750));
  jand g0109(.dina(n750), .dinb(\in2[8] ), .dout(n751));
  jnot g0110(.din(\in2[8] ), .dout(n752));
  jand g0111(.dina(\in3[8] ), .dinb(n752), .dout(n753));
  jnot g0112(.din(n753), .dout(n754));
  jnot g0113(.din(\in3[7] ), .dout(n755));
  jand g0114(.dina(n755), .dinb(\in2[7] ), .dout(n756));
  jnot g0115(.din(\in2[7] ), .dout(n757));
  jand g0116(.dina(\in3[7] ), .dinb(n757), .dout(n758));
  jnot g0117(.din(n758), .dout(n759));
  jnot g0118(.din(\in3[6] ), .dout(n760));
  jand g0119(.dina(n760), .dinb(\in2[6] ), .dout(n761));
  jnot g0120(.din(\in2[6] ), .dout(n762));
  jand g0121(.dina(\in3[6] ), .dinb(n762), .dout(n763));
  jnot g0122(.din(n763), .dout(n764));
  jnot g0123(.din(\in3[5] ), .dout(n765));
  jand g0124(.dina(n765), .dinb(\in2[5] ), .dout(n766));
  jnot g0125(.din(\in2[5] ), .dout(n767));
  jand g0126(.dina(\in3[5] ), .dinb(n767), .dout(n768));
  jnot g0127(.din(n768), .dout(n769));
  jnot g0128(.din(\in3[4] ), .dout(n770));
  jand g0129(.dina(n770), .dinb(\in2[4] ), .dout(n771));
  jnot g0130(.din(\in2[4] ), .dout(n772));
  jand g0131(.dina(\in3[4] ), .dinb(n772), .dout(n773));
  jnot g0132(.din(n773), .dout(n774));
  jnot g0133(.din(\in3[3] ), .dout(n775));
  jand g0134(.dina(n775), .dinb(\in2[3] ), .dout(n776));
  jnot g0135(.din(\in2[3] ), .dout(n777));
  jand g0136(.dina(\in3[3] ), .dinb(n777), .dout(n778));
  jnot g0137(.din(n778), .dout(n779));
  jnot g0138(.din(\in3[2] ), .dout(n780));
  jand g0139(.dina(n780), .dinb(\in2[2] ), .dout(n781));
  jnot g0140(.din(\in2[2] ), .dout(n782));
  jand g0141(.dina(\in3[2] ), .dinb(n782), .dout(n783));
  jnot g0142(.din(n783), .dout(n784));
  jnot g0143(.din(\in3[1] ), .dout(n785));
  jand g0144(.dina(n785), .dinb(\in2[1] ), .dout(n786));
  jor  g0145(.dina(n785), .dinb(\in2[1] ), .dout(n787));
  jnot g0146(.din(\in3[0] ), .dout(n788));
  jand g0147(.dina(n788), .dinb(\in2[0] ), .dout(n789));
  jand g0148(.dina(n789), .dinb(n787), .dout(n790));
  jor  g0149(.dina(n790), .dinb(n786), .dout(n791));
  jand g0150(.dina(n791), .dinb(n784), .dout(n792));
  jor  g0151(.dina(n792), .dinb(n781), .dout(n793));
  jand g0152(.dina(n793), .dinb(n779), .dout(n794));
  jor  g0153(.dina(n794), .dinb(n776), .dout(n795));
  jand g0154(.dina(n795), .dinb(n774), .dout(n796));
  jor  g0155(.dina(n796), .dinb(n771), .dout(n797));
  jand g0156(.dina(n797), .dinb(n769), .dout(n798));
  jor  g0157(.dina(n798), .dinb(n766), .dout(n799));
  jand g0158(.dina(n799), .dinb(n764), .dout(n800));
  jor  g0159(.dina(n800), .dinb(n761), .dout(n801));
  jand g0160(.dina(n801), .dinb(n759), .dout(n802));
  jor  g0161(.dina(n802), .dinb(n756), .dout(n803));
  jand g0162(.dina(n803), .dinb(n754), .dout(n804));
  jor  g0163(.dina(n804), .dinb(n751), .dout(n805));
  jand g0164(.dina(n805), .dinb(n749), .dout(n806));
  jor  g0165(.dina(n806), .dinb(n746), .dout(n807));
  jand g0166(.dina(n807), .dinb(n744), .dout(n808));
  jor  g0167(.dina(n808), .dinb(n741), .dout(n809));
  jand g0168(.dina(n809), .dinb(n739), .dout(n810));
  jor  g0169(.dina(n810), .dinb(n736), .dout(n811));
  jand g0170(.dina(n811), .dinb(n734), .dout(n812));
  jor  g0171(.dina(n812), .dinb(n731), .dout(n813));
  jand g0172(.dina(n813), .dinb(n729), .dout(n814));
  jor  g0173(.dina(n814), .dinb(n726), .dout(n815));
  jand g0174(.dina(n815), .dinb(n724), .dout(n816));
  jor  g0175(.dina(n816), .dinb(n721), .dout(n817));
  jand g0176(.dina(n817), .dinb(n719), .dout(n818));
  jor  g0177(.dina(n818), .dinb(n716), .dout(n819));
  jand g0178(.dina(n819), .dinb(n714), .dout(n820));
  jor  g0179(.dina(n820), .dinb(n711), .dout(n821));
  jand g0180(.dina(n821), .dinb(n709), .dout(n822));
  jor  g0181(.dina(n822), .dinb(n706), .dout(n823));
  jand g0182(.dina(n823), .dinb(n704), .dout(n824));
  jor  g0183(.dina(n824), .dinb(n701), .dout(n825));
  jand g0184(.dina(n825), .dinb(n699), .dout(n826));
  jor  g0185(.dina(n826), .dinb(n696), .dout(n827));
  jand g0186(.dina(n827), .dinb(n694), .dout(n828));
  jor  g0187(.dina(n828), .dinb(n691), .dout(n829));
  jand g0188(.dina(n829), .dinb(n689), .dout(n830));
  jor  g0189(.dina(n830), .dinb(n686), .dout(n831));
  jand g0190(.dina(n831), .dinb(n684), .dout(n832));
  jor  g0191(.dina(n832), .dinb(n681), .dout(n833));
  jand g0192(.dina(n833), .dinb(n679), .dout(n834));
  jor  g0193(.dina(n834), .dinb(n676), .dout(n835));
  jand g0194(.dina(n835), .dinb(n674), .dout(n836));
  jor  g0195(.dina(n836), .dinb(n671), .dout(n837));
  jand g0196(.dina(n837), .dinb(n669), .dout(n838));
  jor  g0197(.dina(n838), .dinb(n666), .dout(n839));
  jand g0198(.dina(n839), .dinb(n664), .dout(n840));
  jor  g0199(.dina(n840), .dinb(n661), .dout(n841));
  jand g0200(.dina(n841), .dinb(n659), .dout(n842));
  jor  g0201(.dina(n842), .dinb(n656), .dout(n843));
  jand g0202(.dina(n843), .dinb(n654), .dout(n844));
  jor  g0203(.dina(n844), .dinb(n651), .dout(n845));
  jand g0204(.dina(n845), .dinb(n649), .dout(n846));
  jor  g0205(.dina(n846), .dinb(n646), .dout(n847));
  jand g0206(.dina(n847), .dinb(n644), .dout(n848));
  jnot g0207(.din(\in3[30] ), .dout(n849));
  jand g0208(.dina(n849), .dinb(\in2[30] ), .dout(n850));
  jnot g0209(.din(\in3[31] ), .dout(n851));
  jand g0210(.dina(n851), .dinb(\in2[31] ), .dout(n852));
  jor  g0211(.dina(n852), .dinb(n850), .dout(n853));
  jor  g0212(.dina(n853), .dinb(n848), .dout(n854));
  jnot g0213(.din(\in2[37] ), .dout(n855));
  jand g0214(.dina(\in3[37] ), .dinb(n855), .dout(n856));
  jnot g0215(.din(\in2[39] ), .dout(n857));
  jand g0216(.dina(\in3[39] ), .dinb(n857), .dout(n858));
  jnot g0217(.din(\in2[38] ), .dout(n859));
  jand g0218(.dina(\in3[38] ), .dinb(n859), .dout(n860));
  jor  g0219(.dina(n860), .dinb(n858), .dout(n861));
  jor  g0220(.dina(n861), .dinb(n856), .dout(n862));
  jnot g0221(.din(\in2[35] ), .dout(n863));
  jand g0222(.dina(\in3[35] ), .dinb(n863), .dout(n864));
  jnot g0223(.din(\in2[34] ), .dout(n865));
  jand g0224(.dina(\in3[34] ), .dinb(n865), .dout(n866));
  jor  g0225(.dina(n866), .dinb(n864), .dout(n867));
  jnot g0226(.din(\in2[32] ), .dout(n868));
  jand g0227(.dina(\in3[32] ), .dinb(n868), .dout(n869));
  jnot g0228(.din(\in2[33] ), .dout(n870));
  jand g0229(.dina(\in3[33] ), .dinb(n870), .dout(n871));
  jor  g0230(.dina(n871), .dinb(n869), .dout(n872));
  jnot g0231(.din(\in2[36] ), .dout(n873));
  jand g0232(.dina(\in3[36] ), .dinb(n873), .dout(n874));
  jnot g0233(.din(\in2[31] ), .dout(n875));
  jand g0234(.dina(\in3[31] ), .dinb(n875), .dout(n876));
  jor  g0235(.dina(n876), .dinb(n874), .dout(n877));
  jor  g0236(.dina(n877), .dinb(n872), .dout(n878));
  jor  g0237(.dina(n878), .dinb(n867), .dout(n879));
  jor  g0238(.dina(n879), .dinb(n862), .dout(n880));
  jnot g0239(.din(n880), .dout(n881));
  jand g0240(.dina(n881), .dinb(n854), .dout(n882));
  jnot g0241(.din(n862), .dout(n883));
  jnot g0242(.din(n874), .dout(n884));
  jnot g0243(.din(\in3[35] ), .dout(n885));
  jand g0244(.dina(n885), .dinb(\in2[35] ), .dout(n886));
  jnot g0245(.din(n867), .dout(n887));
  jnot g0246(.din(n871), .dout(n888));
  jnot g0247(.din(\in3[32] ), .dout(n889));
  jand g0248(.dina(n889), .dinb(\in2[32] ), .dout(n890));
  jand g0249(.dina(n890), .dinb(n888), .dout(n891));
  jnot g0250(.din(\in3[33] ), .dout(n892));
  jand g0251(.dina(n892), .dinb(\in2[33] ), .dout(n893));
  jnot g0252(.din(\in3[34] ), .dout(n894));
  jand g0253(.dina(n894), .dinb(\in2[34] ), .dout(n895));
  jor  g0254(.dina(n895), .dinb(n893), .dout(n896));
  jor  g0255(.dina(n896), .dinb(n891), .dout(n897));
  jand g0256(.dina(n897), .dinb(n887), .dout(n898));
  jor  g0257(.dina(n898), .dinb(n886), .dout(n899));
  jand g0258(.dina(n899), .dinb(n884), .dout(n900));
  jnot g0259(.din(\in3[36] ), .dout(n901));
  jand g0260(.dina(n901), .dinb(\in2[36] ), .dout(n902));
  jnot g0261(.din(\in3[37] ), .dout(n903));
  jand g0262(.dina(n903), .dinb(\in2[37] ), .dout(n904));
  jor  g0263(.dina(n904), .dinb(n902), .dout(n905));
  jor  g0264(.dina(n905), .dinb(n900), .dout(n906));
  jand g0265(.dina(n906), .dinb(n883), .dout(n907));
  jnot g0266(.din(n858), .dout(n908));
  jnot g0267(.din(\in3[38] ), .dout(n909));
  jand g0268(.dina(n909), .dinb(\in2[38] ), .dout(n910));
  jand g0269(.dina(n910), .dinb(n908), .dout(n911));
  jnot g0270(.din(\in3[39] ), .dout(n912));
  jand g0271(.dina(n912), .dinb(\in2[39] ), .dout(n913));
  jor  g0272(.dina(n913), .dinb(n911), .dout(n914));
  jor  g0273(.dina(n914), .dinb(n907), .dout(n915));
  jor  g0274(.dina(n915), .dinb(n882), .dout(n916));
  jnot g0275(.din(\in2[45] ), .dout(n917));
  jand g0276(.dina(\in3[45] ), .dinb(n917), .dout(n918));
  jnot g0277(.din(\in2[47] ), .dout(n919));
  jand g0278(.dina(\in3[47] ), .dinb(n919), .dout(n920));
  jnot g0279(.din(\in2[46] ), .dout(n921));
  jand g0280(.dina(\in3[46] ), .dinb(n921), .dout(n922));
  jor  g0281(.dina(n922), .dinb(n920), .dout(n923));
  jor  g0282(.dina(n923), .dinb(n918), .dout(n924));
  jnot g0283(.din(\in2[43] ), .dout(n925));
  jand g0284(.dina(\in3[43] ), .dinb(n925), .dout(n926));
  jnot g0285(.din(\in2[42] ), .dout(n927));
  jand g0286(.dina(\in3[42] ), .dinb(n927), .dout(n928));
  jor  g0287(.dina(n928), .dinb(n926), .dout(n929));
  jnot g0288(.din(\in2[44] ), .dout(n930));
  jand g0289(.dina(\in3[44] ), .dinb(n930), .dout(n931));
  jnot g0290(.din(\in2[40] ), .dout(n932));
  jand g0291(.dina(\in3[40] ), .dinb(n932), .dout(n933));
  jnot g0292(.din(\in2[41] ), .dout(n934));
  jand g0293(.dina(\in3[41] ), .dinb(n934), .dout(n935));
  jor  g0294(.dina(n935), .dinb(n933), .dout(n936));
  jor  g0295(.dina(n936), .dinb(n931), .dout(n937));
  jor  g0296(.dina(n937), .dinb(n929), .dout(n938));
  jor  g0297(.dina(n938), .dinb(n924), .dout(n939));
  jnot g0298(.din(n939), .dout(n940));
  jand g0299(.dina(n940), .dinb(n916), .dout(n941));
  jnot g0300(.din(n924), .dout(n942));
  jnot g0301(.din(n931), .dout(n943));
  jnot g0302(.din(\in3[43] ), .dout(n944));
  jand g0303(.dina(n944), .dinb(\in2[43] ), .dout(n945));
  jnot g0304(.din(n929), .dout(n946));
  jnot g0305(.din(n935), .dout(n947));
  jnot g0306(.din(\in3[40] ), .dout(n948));
  jand g0307(.dina(n948), .dinb(\in2[40] ), .dout(n949));
  jand g0308(.dina(n949), .dinb(n947), .dout(n950));
  jnot g0309(.din(\in3[41] ), .dout(n951));
  jand g0310(.dina(n951), .dinb(\in2[41] ), .dout(n952));
  jnot g0311(.din(\in3[42] ), .dout(n953));
  jand g0312(.dina(n953), .dinb(\in2[42] ), .dout(n954));
  jor  g0313(.dina(n954), .dinb(n952), .dout(n955));
  jor  g0314(.dina(n955), .dinb(n950), .dout(n956));
  jand g0315(.dina(n956), .dinb(n946), .dout(n957));
  jor  g0316(.dina(n957), .dinb(n945), .dout(n958));
  jand g0317(.dina(n958), .dinb(n943), .dout(n959));
  jnot g0318(.din(\in3[44] ), .dout(n960));
  jand g0319(.dina(n960), .dinb(\in2[44] ), .dout(n961));
  jnot g0320(.din(\in3[45] ), .dout(n962));
  jand g0321(.dina(n962), .dinb(\in2[45] ), .dout(n963));
  jor  g0322(.dina(n963), .dinb(n961), .dout(n964));
  jor  g0323(.dina(n964), .dinb(n959), .dout(n965));
  jand g0324(.dina(n965), .dinb(n942), .dout(n966));
  jnot g0325(.din(n920), .dout(n967));
  jnot g0326(.din(\in3[46] ), .dout(n968));
  jand g0327(.dina(n968), .dinb(\in2[46] ), .dout(n969));
  jand g0328(.dina(n969), .dinb(n967), .dout(n970));
  jnot g0329(.din(\in3[47] ), .dout(n971));
  jand g0330(.dina(n971), .dinb(\in2[47] ), .dout(n972));
  jor  g0331(.dina(n972), .dinb(n970), .dout(n973));
  jor  g0332(.dina(n973), .dinb(n966), .dout(n974));
  jor  g0333(.dina(n974), .dinb(n941), .dout(n975));
  jnot g0334(.din(\in3[52] ), .dout(n976));
  jnot g0335(.din(\in2[53] ), .dout(n977));
  jand g0336(.dina(\in3[53] ), .dinb(n977), .dout(n978));
  jnot g0337(.din(n978), .dout(n979));
  jand g0338(.dina(n979), .dinb(n976), .dout(n980));
  jand g0339(.dina(n979), .dinb(\in2[52] ), .dout(n981));
  jor  g0340(.dina(n981), .dinb(n980), .dout(n982));
  jnot g0341(.din(n982), .dout(n983));
  jnot g0342(.din(\in2[55] ), .dout(n984));
  jand g0343(.dina(\in3[55] ), .dinb(n984), .dout(n985));
  jnot g0344(.din(\in2[54] ), .dout(n986));
  jand g0345(.dina(\in3[54] ), .dinb(n986), .dout(n987));
  jor  g0346(.dina(n987), .dinb(n985), .dout(n988));
  jnot g0347(.din(\in2[51] ), .dout(n989));
  jand g0348(.dina(\in3[51] ), .dinb(n989), .dout(n990));
  jnot g0349(.din(\in2[50] ), .dout(n991));
  jand g0350(.dina(\in3[50] ), .dinb(n991), .dout(n992));
  jor  g0351(.dina(n992), .dinb(n990), .dout(n993));
  jnot g0352(.din(\in2[48] ), .dout(n994));
  jand g0353(.dina(\in3[48] ), .dinb(n994), .dout(n995));
  jnot g0354(.din(\in2[49] ), .dout(n996));
  jand g0355(.dina(\in3[49] ), .dinb(n996), .dout(n997));
  jor  g0356(.dina(n997), .dinb(n995), .dout(n998));
  jor  g0357(.dina(n998), .dinb(n993), .dout(n999));
  jor  g0358(.dina(n999), .dinb(n988), .dout(n1000));
  jor  g0359(.dina(n1000), .dinb(n983), .dout(n1001));
  jnot g0360(.din(n1001), .dout(n1002));
  jand g0361(.dina(n1002), .dinb(n975), .dout(n1003));
  jnot g0362(.din(\in3[55] ), .dout(n1004));
  jand g0363(.dina(n1004), .dinb(\in2[55] ), .dout(n1005));
  jnot g0364(.din(n988), .dout(n1006));
  jnot g0365(.din(\in3[51] ), .dout(n1007));
  jand g0366(.dina(n1007), .dinb(\in2[51] ), .dout(n1008));
  jnot g0367(.din(n993), .dout(n1009));
  jnot g0368(.din(n997), .dout(n1010));
  jnot g0369(.din(\in3[48] ), .dout(n1011));
  jand g0370(.dina(n1011), .dinb(\in2[48] ), .dout(n1012));
  jand g0371(.dina(n1012), .dinb(n1010), .dout(n1013));
  jnot g0372(.din(\in3[49] ), .dout(n1014));
  jand g0373(.dina(n1014), .dinb(\in2[49] ), .dout(n1015));
  jnot g0374(.din(\in3[50] ), .dout(n1016));
  jand g0375(.dina(n1016), .dinb(\in2[50] ), .dout(n1017));
  jor  g0376(.dina(n1017), .dinb(n1015), .dout(n1018));
  jor  g0377(.dina(n1018), .dinb(n1013), .dout(n1019));
  jand g0378(.dina(n1019), .dinb(n1009), .dout(n1020));
  jor  g0379(.dina(n1020), .dinb(n1008), .dout(n1021));
  jand g0380(.dina(n1021), .dinb(n982), .dout(n1022));
  jand g0381(.dina(n980), .dinb(\in2[52] ), .dout(n1023));
  jnot g0382(.din(\in3[53] ), .dout(n1024));
  jand g0383(.dina(n1024), .dinb(\in2[53] ), .dout(n1025));
  jnot g0384(.din(\in3[54] ), .dout(n1026));
  jand g0385(.dina(n1026), .dinb(\in2[54] ), .dout(n1027));
  jor  g0386(.dina(n1027), .dinb(n1025), .dout(n1028));
  jor  g0387(.dina(n1028), .dinb(n1023), .dout(n1029));
  jor  g0388(.dina(n1029), .dinb(n1022), .dout(n1030));
  jand g0389(.dina(n1030), .dinb(n1006), .dout(n1031));
  jor  g0390(.dina(n1031), .dinb(n1005), .dout(n1032));
  jor  g0391(.dina(n1032), .dinb(n1003), .dout(n1033));
  jnot g0392(.din(\in2[61] ), .dout(n1034));
  jand g0393(.dina(\in3[61] ), .dinb(n1034), .dout(n1035));
  jnot g0394(.din(\in2[63] ), .dout(n1036));
  jand g0395(.dina(\in3[63] ), .dinb(n1036), .dout(n1037));
  jnot g0396(.din(\in2[62] ), .dout(n1038));
  jand g0397(.dina(\in3[62] ), .dinb(n1038), .dout(n1039));
  jor  g0398(.dina(n1039), .dinb(n1037), .dout(n1040));
  jor  g0399(.dina(n1040), .dinb(n1035), .dout(n1041));
  jnot g0400(.din(\in2[59] ), .dout(n1042));
  jand g0401(.dina(\in3[59] ), .dinb(n1042), .dout(n1043));
  jnot g0402(.din(\in2[58] ), .dout(n1044));
  jand g0403(.dina(\in3[58] ), .dinb(n1044), .dout(n1045));
  jor  g0404(.dina(n1045), .dinb(n1043), .dout(n1046));
  jnot g0405(.din(\in2[60] ), .dout(n1047));
  jand g0406(.dina(\in3[60] ), .dinb(n1047), .dout(n1048));
  jnot g0407(.din(\in2[56] ), .dout(n1049));
  jand g0408(.dina(\in3[56] ), .dinb(n1049), .dout(n1050));
  jnot g0409(.din(\in2[57] ), .dout(n1051));
  jand g0410(.dina(\in3[57] ), .dinb(n1051), .dout(n1052));
  jor  g0411(.dina(n1052), .dinb(n1050), .dout(n1053));
  jor  g0412(.dina(n1053), .dinb(n1048), .dout(n1054));
  jor  g0413(.dina(n1054), .dinb(n1046), .dout(n1055));
  jor  g0414(.dina(n1055), .dinb(n1041), .dout(n1056));
  jnot g0415(.din(n1056), .dout(n1057));
  jand g0416(.dina(n1057), .dinb(n1033), .dout(n1058));
  jnot g0417(.din(n1041), .dout(n1059));
  jnot g0418(.din(n1048), .dout(n1060));
  jnot g0419(.din(\in3[59] ), .dout(n1061));
  jand g0420(.dina(n1061), .dinb(\in2[59] ), .dout(n1062));
  jnot g0421(.din(n1046), .dout(n1063));
  jnot g0422(.din(n1052), .dout(n1064));
  jnot g0423(.din(\in3[56] ), .dout(n1065));
  jand g0424(.dina(n1065), .dinb(\in2[56] ), .dout(n1066));
  jand g0425(.dina(n1066), .dinb(n1064), .dout(n1067));
  jnot g0426(.din(\in3[57] ), .dout(n1068));
  jand g0427(.dina(n1068), .dinb(\in2[57] ), .dout(n1069));
  jnot g0428(.din(\in3[58] ), .dout(n1070));
  jand g0429(.dina(n1070), .dinb(\in2[58] ), .dout(n1071));
  jor  g0430(.dina(n1071), .dinb(n1069), .dout(n1072));
  jor  g0431(.dina(n1072), .dinb(n1067), .dout(n1073));
  jand g0432(.dina(n1073), .dinb(n1063), .dout(n1074));
  jor  g0433(.dina(n1074), .dinb(n1062), .dout(n1075));
  jand g0434(.dina(n1075), .dinb(n1060), .dout(n1076));
  jnot g0435(.din(\in3[60] ), .dout(n1077));
  jand g0436(.dina(n1077), .dinb(\in2[60] ), .dout(n1078));
  jnot g0437(.din(\in3[61] ), .dout(n1079));
  jand g0438(.dina(n1079), .dinb(\in2[61] ), .dout(n1080));
  jor  g0439(.dina(n1080), .dinb(n1078), .dout(n1081));
  jor  g0440(.dina(n1081), .dinb(n1076), .dout(n1082));
  jand g0441(.dina(n1082), .dinb(n1059), .dout(n1083));
  jnot g0442(.din(n1037), .dout(n1084));
  jnot g0443(.din(\in3[62] ), .dout(n1085));
  jand g0444(.dina(n1085), .dinb(\in2[62] ), .dout(n1086));
  jand g0445(.dina(n1086), .dinb(n1084), .dout(n1087));
  jnot g0446(.din(\in3[63] ), .dout(n1088));
  jand g0447(.dina(n1088), .dinb(\in2[63] ), .dout(n1089));
  jor  g0448(.dina(n1089), .dinb(n1087), .dout(n1090));
  jor  g0449(.dina(n1090), .dinb(n1083), .dout(n1091));
  jor  g0450(.dina(n1091), .dinb(n1058), .dout(n1092));
  jnot g0451(.din(\in2[67] ), .dout(n1093));
  jand g0452(.dina(\in3[67] ), .dinb(n1093), .dout(n1094));
  jnot g0453(.din(\in2[66] ), .dout(n1095));
  jand g0454(.dina(\in3[66] ), .dinb(n1095), .dout(n1096));
  jor  g0455(.dina(n1096), .dinb(n1094), .dout(n1097));
  jnot g0456(.din(\in2[65] ), .dout(n1098));
  jand g0457(.dina(\in3[65] ), .dinb(n1098), .dout(n1099));
  jnot g0458(.din(\in2[64] ), .dout(n1100));
  jand g0459(.dina(\in3[64] ), .dinb(n1100), .dout(n1101));
  jor  g0460(.dina(n1101), .dinb(n1099), .dout(n1102));
  jor  g0461(.dina(n1102), .dinb(n1097), .dout(n1103));
  jnot g0462(.din(n1103), .dout(n1104));
  jand g0463(.dina(n1104), .dinb(n1092), .dout(n1105));
  jnot g0464(.din(\in3[67] ), .dout(n1106));
  jand g0465(.dina(n1106), .dinb(\in2[67] ), .dout(n1107));
  jnot g0466(.din(n1097), .dout(n1108));
  jnot g0467(.din(n1099), .dout(n1109));
  jnot g0468(.din(\in3[64] ), .dout(n1110));
  jand g0469(.dina(n1110), .dinb(\in2[64] ), .dout(n1111));
  jand g0470(.dina(n1111), .dinb(n1109), .dout(n1112));
  jnot g0471(.din(\in3[65] ), .dout(n1113));
  jand g0472(.dina(n1113), .dinb(\in2[65] ), .dout(n1114));
  jnot g0473(.din(\in3[66] ), .dout(n1115));
  jand g0474(.dina(n1115), .dinb(\in2[66] ), .dout(n1116));
  jor  g0475(.dina(n1116), .dinb(n1114), .dout(n1117));
  jor  g0476(.dina(n1117), .dinb(n1112), .dout(n1118));
  jand g0477(.dina(n1118), .dinb(n1108), .dout(n1119));
  jor  g0478(.dina(n1119), .dinb(n1107), .dout(n1120));
  jor  g0479(.dina(n1120), .dinb(n1105), .dout(n1121));
  jnot g0480(.din(\in2[68] ), .dout(n1122));
  jand g0481(.dina(\in3[68] ), .dinb(n1122), .dout(n1123));
  jnot g0482(.din(\in2[69] ), .dout(n1124));
  jand g0483(.dina(\in3[69] ), .dinb(n1124), .dout(n1125));
  jnot g0484(.din(\in2[71] ), .dout(n1126));
  jand g0485(.dina(\in3[71] ), .dinb(n1126), .dout(n1127));
  jnot g0486(.din(\in2[70] ), .dout(n1128));
  jand g0487(.dina(\in3[70] ), .dinb(n1128), .dout(n1129));
  jor  g0488(.dina(n1129), .dinb(n1127), .dout(n1130));
  jor  g0489(.dina(n1130), .dinb(n1125), .dout(n1131));
  jor  g0490(.dina(n1131), .dinb(n1123), .dout(n1132));
  jnot g0491(.din(n1132), .dout(n1133));
  jand g0492(.dina(n1133), .dinb(n1121), .dout(n1134));
  jnot g0493(.din(n1131), .dout(n1135));
  jnot g0494(.din(\in3[69] ), .dout(n1136));
  jand g0495(.dina(n1136), .dinb(\in2[69] ), .dout(n1137));
  jnot g0496(.din(\in3[68] ), .dout(n1138));
  jand g0497(.dina(n1138), .dinb(\in2[68] ), .dout(n1139));
  jor  g0498(.dina(n1139), .dinb(n1137), .dout(n1140));
  jand g0499(.dina(n1140), .dinb(n1135), .dout(n1141));
  jnot g0500(.din(\in3[71] ), .dout(n1142));
  jand g0501(.dina(n1142), .dinb(\in2[71] ), .dout(n1143));
  jnot g0502(.din(n1127), .dout(n1144));
  jnot g0503(.din(\in3[70] ), .dout(n1145));
  jand g0504(.dina(n1145), .dinb(\in2[70] ), .dout(n1146));
  jand g0505(.dina(n1146), .dinb(n1144), .dout(n1147));
  jor  g0506(.dina(n1147), .dinb(n1143), .dout(n1148));
  jor  g0507(.dina(n1148), .dinb(n1141), .dout(n1149));
  jor  g0508(.dina(n1149), .dinb(n1134), .dout(n1150));
  jnot g0509(.din(\in2[75] ), .dout(n1151));
  jand g0510(.dina(\in3[75] ), .dinb(n1151), .dout(n1152));
  jnot g0511(.din(\in2[74] ), .dout(n1153));
  jand g0512(.dina(\in3[74] ), .dinb(n1153), .dout(n1154));
  jor  g0513(.dina(n1154), .dinb(n1152), .dout(n1155));
  jnot g0514(.din(\in2[73] ), .dout(n1156));
  jand g0515(.dina(\in3[73] ), .dinb(n1156), .dout(n1157));
  jnot g0516(.din(\in2[72] ), .dout(n1158));
  jand g0517(.dina(\in3[72] ), .dinb(n1158), .dout(n1159));
  jor  g0518(.dina(n1159), .dinb(n1157), .dout(n1160));
  jor  g0519(.dina(n1160), .dinb(n1155), .dout(n1161));
  jnot g0520(.din(n1161), .dout(n1162));
  jand g0521(.dina(n1162), .dinb(n1150), .dout(n1163));
  jnot g0522(.din(\in3[75] ), .dout(n1164));
  jand g0523(.dina(n1164), .dinb(\in2[75] ), .dout(n1165));
  jnot g0524(.din(n1155), .dout(n1166));
  jnot g0525(.din(n1157), .dout(n1167));
  jnot g0526(.din(\in3[72] ), .dout(n1168));
  jand g0527(.dina(n1168), .dinb(\in2[72] ), .dout(n1169));
  jand g0528(.dina(n1169), .dinb(n1167), .dout(n1170));
  jnot g0529(.din(\in3[73] ), .dout(n1171));
  jand g0530(.dina(n1171), .dinb(\in2[73] ), .dout(n1172));
  jnot g0531(.din(\in3[74] ), .dout(n1173));
  jand g0532(.dina(n1173), .dinb(\in2[74] ), .dout(n1174));
  jor  g0533(.dina(n1174), .dinb(n1172), .dout(n1175));
  jor  g0534(.dina(n1175), .dinb(n1170), .dout(n1176));
  jand g0535(.dina(n1176), .dinb(n1166), .dout(n1177));
  jor  g0536(.dina(n1177), .dinb(n1165), .dout(n1178));
  jor  g0537(.dina(n1178), .dinb(n1163), .dout(n1179));
  jnot g0538(.din(\in2[76] ), .dout(n1180));
  jand g0539(.dina(\in3[76] ), .dinb(n1180), .dout(n1181));
  jnot g0540(.din(\in2[77] ), .dout(n1182));
  jand g0541(.dina(\in3[77] ), .dinb(n1182), .dout(n1183));
  jnot g0542(.din(\in2[79] ), .dout(n1184));
  jand g0543(.dina(\in3[79] ), .dinb(n1184), .dout(n1185));
  jnot g0544(.din(\in2[78] ), .dout(n1186));
  jand g0545(.dina(\in3[78] ), .dinb(n1186), .dout(n1187));
  jor  g0546(.dina(n1187), .dinb(n1185), .dout(n1188));
  jor  g0547(.dina(n1188), .dinb(n1183), .dout(n1189));
  jor  g0548(.dina(n1189), .dinb(n1181), .dout(n1190));
  jnot g0549(.din(n1190), .dout(n1191));
  jand g0550(.dina(n1191), .dinb(n1179), .dout(n1192));
  jnot g0551(.din(n1189), .dout(n1193));
  jnot g0552(.din(\in3[77] ), .dout(n1194));
  jand g0553(.dina(n1194), .dinb(\in2[77] ), .dout(n1195));
  jnot g0554(.din(\in3[76] ), .dout(n1196));
  jand g0555(.dina(n1196), .dinb(\in2[76] ), .dout(n1197));
  jor  g0556(.dina(n1197), .dinb(n1195), .dout(n1198));
  jand g0557(.dina(n1198), .dinb(n1193), .dout(n1199));
  jnot g0558(.din(\in3[79] ), .dout(n1200));
  jand g0559(.dina(n1200), .dinb(\in2[79] ), .dout(n1201));
  jnot g0560(.din(n1185), .dout(n1202));
  jnot g0561(.din(\in3[78] ), .dout(n1203));
  jand g0562(.dina(n1203), .dinb(\in2[78] ), .dout(n1204));
  jand g0563(.dina(n1204), .dinb(n1202), .dout(n1205));
  jor  g0564(.dina(n1205), .dinb(n1201), .dout(n1206));
  jor  g0565(.dina(n1206), .dinb(n1199), .dout(n1207));
  jor  g0566(.dina(n1207), .dinb(n1192), .dout(n1208));
  jnot g0567(.din(\in2[83] ), .dout(n1209));
  jand g0568(.dina(\in3[83] ), .dinb(n1209), .dout(n1210));
  jnot g0569(.din(\in2[82] ), .dout(n1211));
  jand g0570(.dina(\in3[82] ), .dinb(n1211), .dout(n1212));
  jor  g0571(.dina(n1212), .dinb(n1210), .dout(n1213));
  jnot g0572(.din(\in2[81] ), .dout(n1214));
  jand g0573(.dina(\in3[81] ), .dinb(n1214), .dout(n1215));
  jnot g0574(.din(\in2[80] ), .dout(n1216));
  jand g0575(.dina(\in3[80] ), .dinb(n1216), .dout(n1217));
  jor  g0576(.dina(n1217), .dinb(n1215), .dout(n1218));
  jor  g0577(.dina(n1218), .dinb(n1213), .dout(n1219));
  jnot g0578(.din(n1219), .dout(n1220));
  jand g0579(.dina(n1220), .dinb(n1208), .dout(n1221));
  jnot g0580(.din(\in3[83] ), .dout(n1222));
  jand g0581(.dina(n1222), .dinb(\in2[83] ), .dout(n1223));
  jnot g0582(.din(n1213), .dout(n1224));
  jnot g0583(.din(n1215), .dout(n1225));
  jnot g0584(.din(\in3[80] ), .dout(n1226));
  jand g0585(.dina(n1226), .dinb(\in2[80] ), .dout(n1227));
  jand g0586(.dina(n1227), .dinb(n1225), .dout(n1228));
  jnot g0587(.din(\in3[81] ), .dout(n1229));
  jand g0588(.dina(n1229), .dinb(\in2[81] ), .dout(n1230));
  jnot g0589(.din(\in3[82] ), .dout(n1231));
  jand g0590(.dina(n1231), .dinb(\in2[82] ), .dout(n1232));
  jor  g0591(.dina(n1232), .dinb(n1230), .dout(n1233));
  jor  g0592(.dina(n1233), .dinb(n1228), .dout(n1234));
  jand g0593(.dina(n1234), .dinb(n1224), .dout(n1235));
  jor  g0594(.dina(n1235), .dinb(n1223), .dout(n1236));
  jor  g0595(.dina(n1236), .dinb(n1221), .dout(n1237));
  jnot g0596(.din(\in2[84] ), .dout(n1238));
  jand g0597(.dina(\in3[84] ), .dinb(n1238), .dout(n1239));
  jnot g0598(.din(\in2[85] ), .dout(n1240));
  jand g0599(.dina(\in3[85] ), .dinb(n1240), .dout(n1241));
  jnot g0600(.din(\in2[87] ), .dout(n1242));
  jand g0601(.dina(\in3[87] ), .dinb(n1242), .dout(n1243));
  jnot g0602(.din(\in2[86] ), .dout(n1244));
  jand g0603(.dina(\in3[86] ), .dinb(n1244), .dout(n1245));
  jor  g0604(.dina(n1245), .dinb(n1243), .dout(n1246));
  jor  g0605(.dina(n1246), .dinb(n1241), .dout(n1247));
  jor  g0606(.dina(n1247), .dinb(n1239), .dout(n1248));
  jnot g0607(.din(n1248), .dout(n1249));
  jand g0608(.dina(n1249), .dinb(n1237), .dout(n1250));
  jnot g0609(.din(n1247), .dout(n1251));
  jnot g0610(.din(\in3[85] ), .dout(n1252));
  jand g0611(.dina(n1252), .dinb(\in2[85] ), .dout(n1253));
  jnot g0612(.din(\in3[84] ), .dout(n1254));
  jand g0613(.dina(n1254), .dinb(\in2[84] ), .dout(n1255));
  jor  g0614(.dina(n1255), .dinb(n1253), .dout(n1256));
  jand g0615(.dina(n1256), .dinb(n1251), .dout(n1257));
  jnot g0616(.din(\in3[87] ), .dout(n1258));
  jand g0617(.dina(n1258), .dinb(\in2[87] ), .dout(n1259));
  jnot g0618(.din(n1243), .dout(n1260));
  jnot g0619(.din(\in3[86] ), .dout(n1261));
  jand g0620(.dina(n1261), .dinb(\in2[86] ), .dout(n1262));
  jand g0621(.dina(n1262), .dinb(n1260), .dout(n1263));
  jor  g0622(.dina(n1263), .dinb(n1259), .dout(n1264));
  jor  g0623(.dina(n1264), .dinb(n1257), .dout(n1265));
  jor  g0624(.dina(n1265), .dinb(n1250), .dout(n1266));
  jnot g0625(.din(\in2[91] ), .dout(n1267));
  jand g0626(.dina(\in3[91] ), .dinb(n1267), .dout(n1268));
  jnot g0627(.din(\in2[90] ), .dout(n1269));
  jand g0628(.dina(\in3[90] ), .dinb(n1269), .dout(n1270));
  jor  g0629(.dina(n1270), .dinb(n1268), .dout(n1271));
  jnot g0630(.din(\in2[89] ), .dout(n1272));
  jand g0631(.dina(\in3[89] ), .dinb(n1272), .dout(n1273));
  jnot g0632(.din(\in2[88] ), .dout(n1274));
  jand g0633(.dina(\in3[88] ), .dinb(n1274), .dout(n1275));
  jor  g0634(.dina(n1275), .dinb(n1273), .dout(n1276));
  jor  g0635(.dina(n1276), .dinb(n1271), .dout(n1277));
  jnot g0636(.din(n1277), .dout(n1278));
  jand g0637(.dina(n1278), .dinb(n1266), .dout(n1279));
  jnot g0638(.din(\in3[91] ), .dout(n1280));
  jand g0639(.dina(n1280), .dinb(\in2[91] ), .dout(n1281));
  jnot g0640(.din(n1271), .dout(n1282));
  jnot g0641(.din(n1273), .dout(n1283));
  jnot g0642(.din(\in3[88] ), .dout(n1284));
  jand g0643(.dina(n1284), .dinb(\in2[88] ), .dout(n1285));
  jand g0644(.dina(n1285), .dinb(n1283), .dout(n1286));
  jnot g0645(.din(\in3[89] ), .dout(n1287));
  jand g0646(.dina(n1287), .dinb(\in2[89] ), .dout(n1288));
  jnot g0647(.din(\in3[90] ), .dout(n1289));
  jand g0648(.dina(n1289), .dinb(\in2[90] ), .dout(n1290));
  jor  g0649(.dina(n1290), .dinb(n1288), .dout(n1291));
  jor  g0650(.dina(n1291), .dinb(n1286), .dout(n1292));
  jand g0651(.dina(n1292), .dinb(n1282), .dout(n1293));
  jor  g0652(.dina(n1293), .dinb(n1281), .dout(n1294));
  jor  g0653(.dina(n1294), .dinb(n1279), .dout(n1295));
  jnot g0654(.din(\in2[92] ), .dout(n1296));
  jand g0655(.dina(\in3[92] ), .dinb(n1296), .dout(n1297));
  jnot g0656(.din(\in2[93] ), .dout(n1298));
  jand g0657(.dina(\in3[93] ), .dinb(n1298), .dout(n1299));
  jnot g0658(.din(\in2[95] ), .dout(n1300));
  jand g0659(.dina(\in3[95] ), .dinb(n1300), .dout(n1301));
  jnot g0660(.din(\in2[94] ), .dout(n1302));
  jand g0661(.dina(\in3[94] ), .dinb(n1302), .dout(n1303));
  jor  g0662(.dina(n1303), .dinb(n1301), .dout(n1304));
  jor  g0663(.dina(n1304), .dinb(n1299), .dout(n1305));
  jor  g0664(.dina(n1305), .dinb(n1297), .dout(n1306));
  jnot g0665(.din(n1306), .dout(n1307));
  jand g0666(.dina(n1307), .dinb(n1295), .dout(n1308));
  jnot g0667(.din(n1305), .dout(n1309));
  jnot g0668(.din(\in3[93] ), .dout(n1310));
  jand g0669(.dina(n1310), .dinb(\in2[93] ), .dout(n1311));
  jnot g0670(.din(\in3[92] ), .dout(n1312));
  jand g0671(.dina(n1312), .dinb(\in2[92] ), .dout(n1313));
  jor  g0672(.dina(n1313), .dinb(n1311), .dout(n1314));
  jand g0673(.dina(n1314), .dinb(n1309), .dout(n1315));
  jnot g0674(.din(\in3[95] ), .dout(n1316));
  jand g0675(.dina(n1316), .dinb(\in2[95] ), .dout(n1317));
  jnot g0676(.din(n1301), .dout(n1318));
  jnot g0677(.din(\in3[94] ), .dout(n1319));
  jand g0678(.dina(n1319), .dinb(\in2[94] ), .dout(n1320));
  jand g0679(.dina(n1320), .dinb(n1318), .dout(n1321));
  jor  g0680(.dina(n1321), .dinb(n1317), .dout(n1322));
  jor  g0681(.dina(n1322), .dinb(n1315), .dout(n1323));
  jor  g0682(.dina(n1323), .dinb(n1308), .dout(n1324));
  jnot g0683(.din(\in2[99] ), .dout(n1325));
  jand g0684(.dina(\in3[99] ), .dinb(n1325), .dout(n1326));
  jnot g0685(.din(\in2[98] ), .dout(n1327));
  jand g0686(.dina(\in3[98] ), .dinb(n1327), .dout(n1328));
  jor  g0687(.dina(n1328), .dinb(n1326), .dout(n1329));
  jnot g0688(.din(\in2[97] ), .dout(n1330));
  jand g0689(.dina(\in3[97] ), .dinb(n1330), .dout(n1331));
  jnot g0690(.din(\in2[96] ), .dout(n1332));
  jand g0691(.dina(\in3[96] ), .dinb(n1332), .dout(n1333));
  jor  g0692(.dina(n1333), .dinb(n1331), .dout(n1334));
  jor  g0693(.dina(n1334), .dinb(n1329), .dout(n1335));
  jnot g0694(.din(n1335), .dout(n1336));
  jand g0695(.dina(n1336), .dinb(n1324), .dout(n1337));
  jnot g0696(.din(\in3[99] ), .dout(n1338));
  jand g0697(.dina(n1338), .dinb(\in2[99] ), .dout(n1339));
  jnot g0698(.din(n1329), .dout(n1340));
  jnot g0699(.din(n1331), .dout(n1341));
  jnot g0700(.din(\in3[96] ), .dout(n1342));
  jand g0701(.dina(n1342), .dinb(\in2[96] ), .dout(n1343));
  jand g0702(.dina(n1343), .dinb(n1341), .dout(n1344));
  jnot g0703(.din(\in3[97] ), .dout(n1345));
  jand g0704(.dina(n1345), .dinb(\in2[97] ), .dout(n1346));
  jnot g0705(.din(\in3[98] ), .dout(n1347));
  jand g0706(.dina(n1347), .dinb(\in2[98] ), .dout(n1348));
  jor  g0707(.dina(n1348), .dinb(n1346), .dout(n1349));
  jor  g0708(.dina(n1349), .dinb(n1344), .dout(n1350));
  jand g0709(.dina(n1350), .dinb(n1340), .dout(n1351));
  jor  g0710(.dina(n1351), .dinb(n1339), .dout(n1352));
  jor  g0711(.dina(n1352), .dinb(n1337), .dout(n1353));
  jnot g0712(.din(\in2[100] ), .dout(n1354));
  jand g0713(.dina(\in3[100] ), .dinb(n1354), .dout(n1355));
  jnot g0714(.din(\in2[101] ), .dout(n1356));
  jand g0715(.dina(\in3[101] ), .dinb(n1356), .dout(n1357));
  jnot g0716(.din(\in2[103] ), .dout(n1358));
  jand g0717(.dina(\in3[103] ), .dinb(n1358), .dout(n1359));
  jnot g0718(.din(\in2[102] ), .dout(n1360));
  jand g0719(.dina(\in3[102] ), .dinb(n1360), .dout(n1361));
  jor  g0720(.dina(n1361), .dinb(n1359), .dout(n1362));
  jor  g0721(.dina(n1362), .dinb(n1357), .dout(n1363));
  jor  g0722(.dina(n1363), .dinb(n1355), .dout(n1364));
  jnot g0723(.din(n1364), .dout(n1365));
  jand g0724(.dina(n1365), .dinb(n1353), .dout(n1366));
  jnot g0725(.din(n1363), .dout(n1367));
  jnot g0726(.din(\in3[101] ), .dout(n1368));
  jand g0727(.dina(n1368), .dinb(\in2[101] ), .dout(n1369));
  jnot g0728(.din(\in3[100] ), .dout(n1370));
  jand g0729(.dina(n1370), .dinb(\in2[100] ), .dout(n1371));
  jor  g0730(.dina(n1371), .dinb(n1369), .dout(n1372));
  jand g0731(.dina(n1372), .dinb(n1367), .dout(n1373));
  jnot g0732(.din(\in3[103] ), .dout(n1374));
  jand g0733(.dina(n1374), .dinb(\in2[103] ), .dout(n1375));
  jnot g0734(.din(n1359), .dout(n1376));
  jnot g0735(.din(\in3[102] ), .dout(n1377));
  jand g0736(.dina(n1377), .dinb(\in2[102] ), .dout(n1378));
  jand g0737(.dina(n1378), .dinb(n1376), .dout(n1379));
  jor  g0738(.dina(n1379), .dinb(n1375), .dout(n1380));
  jor  g0739(.dina(n1380), .dinb(n1373), .dout(n1381));
  jor  g0740(.dina(n1381), .dinb(n1366), .dout(n1382));
  jnot g0741(.din(\in2[107] ), .dout(n1383));
  jand g0742(.dina(\in3[107] ), .dinb(n1383), .dout(n1384));
  jnot g0743(.din(\in2[106] ), .dout(n1385));
  jand g0744(.dina(\in3[106] ), .dinb(n1385), .dout(n1386));
  jor  g0745(.dina(n1386), .dinb(n1384), .dout(n1387));
  jnot g0746(.din(\in2[105] ), .dout(n1388));
  jand g0747(.dina(\in3[105] ), .dinb(n1388), .dout(n1389));
  jnot g0748(.din(\in2[104] ), .dout(n1390));
  jand g0749(.dina(\in3[104] ), .dinb(n1390), .dout(n1391));
  jor  g0750(.dina(n1391), .dinb(n1389), .dout(n1392));
  jor  g0751(.dina(n1392), .dinb(n1387), .dout(n1393));
  jnot g0752(.din(n1393), .dout(n1394));
  jand g0753(.dina(n1394), .dinb(n1382), .dout(n1395));
  jnot g0754(.din(\in3[107] ), .dout(n1396));
  jand g0755(.dina(n1396), .dinb(\in2[107] ), .dout(n1397));
  jnot g0756(.din(n1387), .dout(n1398));
  jnot g0757(.din(n1389), .dout(n1399));
  jnot g0758(.din(\in3[104] ), .dout(n1400));
  jand g0759(.dina(n1400), .dinb(\in2[104] ), .dout(n1401));
  jand g0760(.dina(n1401), .dinb(n1399), .dout(n1402));
  jnot g0761(.din(\in3[105] ), .dout(n1403));
  jand g0762(.dina(n1403), .dinb(\in2[105] ), .dout(n1404));
  jnot g0763(.din(\in3[106] ), .dout(n1405));
  jand g0764(.dina(n1405), .dinb(\in2[106] ), .dout(n1406));
  jor  g0765(.dina(n1406), .dinb(n1404), .dout(n1407));
  jor  g0766(.dina(n1407), .dinb(n1402), .dout(n1408));
  jand g0767(.dina(n1408), .dinb(n1398), .dout(n1409));
  jor  g0768(.dina(n1409), .dinb(n1397), .dout(n1410));
  jor  g0769(.dina(n1410), .dinb(n1395), .dout(n1411));
  jnot g0770(.din(\in2[108] ), .dout(n1412));
  jand g0771(.dina(\in3[108] ), .dinb(n1412), .dout(n1413));
  jnot g0772(.din(\in2[109] ), .dout(n1414));
  jand g0773(.dina(\in3[109] ), .dinb(n1414), .dout(n1415));
  jnot g0774(.din(\in2[111] ), .dout(n1416));
  jand g0775(.dina(\in3[111] ), .dinb(n1416), .dout(n1417));
  jnot g0776(.din(\in2[110] ), .dout(n1418));
  jand g0777(.dina(\in3[110] ), .dinb(n1418), .dout(n1419));
  jor  g0778(.dina(n1419), .dinb(n1417), .dout(n1420));
  jor  g0779(.dina(n1420), .dinb(n1415), .dout(n1421));
  jor  g0780(.dina(n1421), .dinb(n1413), .dout(n1422));
  jnot g0781(.din(n1422), .dout(n1423));
  jand g0782(.dina(n1423), .dinb(n1411), .dout(n1424));
  jnot g0783(.din(n1421), .dout(n1425));
  jnot g0784(.din(\in3[109] ), .dout(n1426));
  jand g0785(.dina(n1426), .dinb(\in2[109] ), .dout(n1427));
  jnot g0786(.din(\in3[108] ), .dout(n1428));
  jand g0787(.dina(n1428), .dinb(\in2[108] ), .dout(n1429));
  jor  g0788(.dina(n1429), .dinb(n1427), .dout(n1430));
  jand g0789(.dina(n1430), .dinb(n1425), .dout(n1431));
  jnot g0790(.din(\in3[111] ), .dout(n1432));
  jand g0791(.dina(n1432), .dinb(\in2[111] ), .dout(n1433));
  jnot g0792(.din(n1417), .dout(n1434));
  jnot g0793(.din(\in3[110] ), .dout(n1435));
  jand g0794(.dina(n1435), .dinb(\in2[110] ), .dout(n1436));
  jand g0795(.dina(n1436), .dinb(n1434), .dout(n1437));
  jor  g0796(.dina(n1437), .dinb(n1433), .dout(n1438));
  jor  g0797(.dina(n1438), .dinb(n1431), .dout(n1439));
  jor  g0798(.dina(n1439), .dinb(n1424), .dout(n1440));
  jnot g0799(.din(\in2[115] ), .dout(n1441));
  jand g0800(.dina(\in3[115] ), .dinb(n1441), .dout(n1442));
  jnot g0801(.din(\in2[114] ), .dout(n1443));
  jand g0802(.dina(\in3[114] ), .dinb(n1443), .dout(n1444));
  jor  g0803(.dina(n1444), .dinb(n1442), .dout(n1445));
  jnot g0804(.din(\in2[113] ), .dout(n1446));
  jand g0805(.dina(\in3[113] ), .dinb(n1446), .dout(n1447));
  jnot g0806(.din(\in2[112] ), .dout(n1448));
  jand g0807(.dina(\in3[112] ), .dinb(n1448), .dout(n1449));
  jor  g0808(.dina(n1449), .dinb(n1447), .dout(n1450));
  jor  g0809(.dina(n1450), .dinb(n1445), .dout(n1451));
  jnot g0810(.din(n1451), .dout(n1452));
  jand g0811(.dina(n1452), .dinb(n1440), .dout(n1453));
  jnot g0812(.din(\in3[115] ), .dout(n1454));
  jand g0813(.dina(n1454), .dinb(\in2[115] ), .dout(n1455));
  jnot g0814(.din(n1445), .dout(n1456));
  jnot g0815(.din(n1447), .dout(n1457));
  jnot g0816(.din(\in3[112] ), .dout(n1458));
  jand g0817(.dina(n1458), .dinb(\in2[112] ), .dout(n1459));
  jand g0818(.dina(n1459), .dinb(n1457), .dout(n1460));
  jnot g0819(.din(\in3[113] ), .dout(n1461));
  jand g0820(.dina(n1461), .dinb(\in2[113] ), .dout(n1462));
  jnot g0821(.din(\in3[114] ), .dout(n1463));
  jand g0822(.dina(n1463), .dinb(\in2[114] ), .dout(n1464));
  jor  g0823(.dina(n1464), .dinb(n1462), .dout(n1465));
  jor  g0824(.dina(n1465), .dinb(n1460), .dout(n1466));
  jand g0825(.dina(n1466), .dinb(n1456), .dout(n1467));
  jor  g0826(.dina(n1467), .dinb(n1455), .dout(n1468));
  jor  g0827(.dina(n1468), .dinb(n1453), .dout(n1469));
  jnot g0828(.din(\in2[116] ), .dout(n1470));
  jand g0829(.dina(\in3[116] ), .dinb(n1470), .dout(n1471));
  jnot g0830(.din(\in2[117] ), .dout(n1472));
  jand g0831(.dina(\in3[117] ), .dinb(n1472), .dout(n1473));
  jnot g0832(.din(\in2[119] ), .dout(n1474));
  jand g0833(.dina(\in3[119] ), .dinb(n1474), .dout(n1475));
  jnot g0834(.din(\in2[118] ), .dout(n1476));
  jand g0835(.dina(\in3[118] ), .dinb(n1476), .dout(n1477));
  jor  g0836(.dina(n1477), .dinb(n1475), .dout(n1478));
  jor  g0837(.dina(n1478), .dinb(n1473), .dout(n1479));
  jor  g0838(.dina(n1479), .dinb(n1471), .dout(n1480));
  jnot g0839(.din(n1480), .dout(n1481));
  jand g0840(.dina(n1481), .dinb(n1469), .dout(n1482));
  jnot g0841(.din(n1479), .dout(n1483));
  jnot g0842(.din(\in3[117] ), .dout(n1484));
  jand g0843(.dina(n1484), .dinb(\in2[117] ), .dout(n1485));
  jnot g0844(.din(\in3[116] ), .dout(n1486));
  jand g0845(.dina(n1486), .dinb(\in2[116] ), .dout(n1487));
  jor  g0846(.dina(n1487), .dinb(n1485), .dout(n1488));
  jand g0847(.dina(n1488), .dinb(n1483), .dout(n1489));
  jnot g0848(.din(\in3[119] ), .dout(n1490));
  jand g0849(.dina(n1490), .dinb(\in2[119] ), .dout(n1491));
  jnot g0850(.din(n1475), .dout(n1492));
  jnot g0851(.din(\in3[118] ), .dout(n1493));
  jand g0852(.dina(n1493), .dinb(\in2[118] ), .dout(n1494));
  jand g0853(.dina(n1494), .dinb(n1492), .dout(n1495));
  jor  g0854(.dina(n1495), .dinb(n1491), .dout(n1496));
  jor  g0855(.dina(n1496), .dinb(n1489), .dout(n1497));
  jor  g0856(.dina(n1497), .dinb(n1482), .dout(n1498));
  jnot g0857(.din(\in2[123] ), .dout(n1499));
  jand g0858(.dina(\in3[123] ), .dinb(n1499), .dout(n1500));
  jnot g0859(.din(\in2[122] ), .dout(n1501));
  jand g0860(.dina(\in3[122] ), .dinb(n1501), .dout(n1502));
  jor  g0861(.dina(n1502), .dinb(n1500), .dout(n1503));
  jnot g0862(.din(\in2[121] ), .dout(n1504));
  jand g0863(.dina(\in3[121] ), .dinb(n1504), .dout(n1505));
  jnot g0864(.din(\in2[120] ), .dout(n1506));
  jand g0865(.dina(\in3[120] ), .dinb(n1506), .dout(n1507));
  jor  g0866(.dina(n1507), .dinb(n1505), .dout(n1508));
  jor  g0867(.dina(n1508), .dinb(n1503), .dout(n1509));
  jnot g0868(.din(n1509), .dout(n1510));
  jand g0869(.dina(n1510), .dinb(n1498), .dout(n1511));
  jnot g0870(.din(\in3[123] ), .dout(n1512));
  jand g0871(.dina(n1512), .dinb(\in2[123] ), .dout(n1513));
  jnot g0872(.din(n1503), .dout(n1514));
  jnot g0873(.din(n1505), .dout(n1515));
  jnot g0874(.din(\in3[120] ), .dout(n1516));
  jand g0875(.dina(n1516), .dinb(\in2[120] ), .dout(n1517));
  jand g0876(.dina(n1517), .dinb(n1515), .dout(n1518));
  jnot g0877(.din(\in3[121] ), .dout(n1519));
  jand g0878(.dina(n1519), .dinb(\in2[121] ), .dout(n1520));
  jnot g0879(.din(\in3[122] ), .dout(n1521));
  jand g0880(.dina(n1521), .dinb(\in2[122] ), .dout(n1522));
  jor  g0881(.dina(n1522), .dinb(n1520), .dout(n1523));
  jor  g0882(.dina(n1523), .dinb(n1518), .dout(n1524));
  jand g0883(.dina(n1524), .dinb(n1514), .dout(n1525));
  jor  g0884(.dina(n1525), .dinb(n1513), .dout(n1526));
  jor  g0885(.dina(n1526), .dinb(n1511), .dout(n1527));
  jnot g0886(.din(\in2[126] ), .dout(n1528));
  jand g0887(.dina(\in3[126] ), .dinb(n1528), .dout(n1529));
  jnot g0888(.din(\in2[125] ), .dout(n1530));
  jand g0889(.dina(\in3[125] ), .dinb(n1530), .dout(n1531));
  jor  g0890(.dina(n1531), .dinb(n1529), .dout(n1532));
  jnot g0891(.din(\in3[127] ), .dout(n1533));
  jand g0892(.dina(n1533), .dinb(\in2[127] ), .dout(n1534));
  jnot g0893(.din(\in2[124] ), .dout(n1535));
  jand g0894(.dina(\in3[124] ), .dinb(n1535), .dout(n1536));
  jor  g0895(.dina(n1536), .dinb(n1534), .dout(n1537));
  jor  g0896(.dina(n1537), .dinb(n1532), .dout(n1538));
  jnot g0897(.din(n1538), .dout(n1539));
  jand g0898(.dina(n1539), .dinb(n1527), .dout(n1540));
  jnot g0899(.din(n1534), .dout(n1541));
  jnot g0900(.din(n1532), .dout(n1542));
  jnot g0901(.din(\in3[124] ), .dout(n1543));
  jand g0902(.dina(n1543), .dinb(\in2[124] ), .dout(n1544));
  jnot g0903(.din(\in3[125] ), .dout(n1545));
  jand g0904(.dina(n1545), .dinb(\in2[125] ), .dout(n1546));
  jor  g0905(.dina(n1546), .dinb(n1544), .dout(n1547));
  jand g0906(.dina(n1547), .dinb(n1542), .dout(n1548));
  jnot g0907(.din(\in3[126] ), .dout(n1549));
  jand g0908(.dina(n1549), .dinb(\in2[126] ), .dout(n1550));
  jor  g0909(.dina(n1550), .dinb(n1548), .dout(n1551));
  jand g0910(.dina(n1551), .dinb(n1541), .dout(n1552));
  jnot g0911(.din(\in2[127] ), .dout(n1553));
  jand g0912(.dina(\in3[127] ), .dinb(n1553), .dout(n1554));
  jor  g0913(.dina(n1554), .dinb(n1552), .dout(n1555));
  jor  g0914(.dina(n1555), .dinb(n1540), .dout(n1556));
  jand g0915(.dina(n1556), .dinb(\in2[0] ), .dout(n1557));
  jnot g0916(.din(n646), .dout(n1558));
  jnot g0917(.din(n651), .dout(n1559));
  jnot g0918(.din(n656), .dout(n1560));
  jnot g0919(.din(n661), .dout(n1561));
  jnot g0920(.din(n666), .dout(n1562));
  jnot g0921(.din(n671), .dout(n1563));
  jnot g0922(.din(n676), .dout(n1564));
  jnot g0923(.din(n681), .dout(n1565));
  jnot g0924(.din(n686), .dout(n1566));
  jnot g0925(.din(n691), .dout(n1567));
  jnot g0926(.din(n696), .dout(n1568));
  jnot g0927(.din(n701), .dout(n1569));
  jnot g0928(.din(n706), .dout(n1570));
  jnot g0929(.din(n711), .dout(n1571));
  jnot g0930(.din(n716), .dout(n1572));
  jnot g0931(.din(n721), .dout(n1573));
  jnot g0932(.din(n726), .dout(n1574));
  jnot g0933(.din(n731), .dout(n1575));
  jnot g0934(.din(n736), .dout(n1576));
  jnot g0935(.din(n741), .dout(n1577));
  jnot g0936(.din(n746), .dout(n1578));
  jnot g0937(.din(n751), .dout(n1579));
  jnot g0938(.din(n756), .dout(n1580));
  jnot g0939(.din(n761), .dout(n1581));
  jnot g0940(.din(n766), .dout(n1582));
  jnot g0941(.din(n771), .dout(n1583));
  jnot g0942(.din(n776), .dout(n1584));
  jnot g0943(.din(n781), .dout(n1585));
  jnot g0944(.din(\in2[1] ), .dout(n1586));
  jor  g0945(.dina(\in3[1] ), .dinb(n1586), .dout(n1587));
  jand g0946(.dina(\in3[1] ), .dinb(n1586), .dout(n1588));
  jnot g0947(.din(\in2[0] ), .dout(n1589));
  jor  g0948(.dina(\in3[0] ), .dinb(n1589), .dout(n1590));
  jor  g0949(.dina(n1590), .dinb(n1588), .dout(n1591));
  jand g0950(.dina(n1591), .dinb(n1587), .dout(n1592));
  jor  g0951(.dina(n1592), .dinb(n783), .dout(n1593));
  jand g0952(.dina(n1593), .dinb(n1585), .dout(n1594));
  jor  g0953(.dina(n1594), .dinb(n778), .dout(n1595));
  jand g0954(.dina(n1595), .dinb(n1584), .dout(n1596));
  jor  g0955(.dina(n1596), .dinb(n773), .dout(n1597));
  jand g0956(.dina(n1597), .dinb(n1583), .dout(n1598));
  jor  g0957(.dina(n1598), .dinb(n768), .dout(n1599));
  jand g0958(.dina(n1599), .dinb(n1582), .dout(n1600));
  jor  g0959(.dina(n1600), .dinb(n763), .dout(n1601));
  jand g0960(.dina(n1601), .dinb(n1581), .dout(n1602));
  jor  g0961(.dina(n1602), .dinb(n758), .dout(n1603));
  jand g0962(.dina(n1603), .dinb(n1580), .dout(n1604));
  jor  g0963(.dina(n1604), .dinb(n753), .dout(n1605));
  jand g0964(.dina(n1605), .dinb(n1579), .dout(n1606));
  jor  g0965(.dina(n1606), .dinb(n748), .dout(n1607));
  jand g0966(.dina(n1607), .dinb(n1578), .dout(n1608));
  jor  g0967(.dina(n1608), .dinb(n743), .dout(n1609));
  jand g0968(.dina(n1609), .dinb(n1577), .dout(n1610));
  jor  g0969(.dina(n1610), .dinb(n738), .dout(n1611));
  jand g0970(.dina(n1611), .dinb(n1576), .dout(n1612));
  jor  g0971(.dina(n1612), .dinb(n733), .dout(n1613));
  jand g0972(.dina(n1613), .dinb(n1575), .dout(n1614));
  jor  g0973(.dina(n1614), .dinb(n728), .dout(n1615));
  jand g0974(.dina(n1615), .dinb(n1574), .dout(n1616));
  jor  g0975(.dina(n1616), .dinb(n723), .dout(n1617));
  jand g0976(.dina(n1617), .dinb(n1573), .dout(n1618));
  jor  g0977(.dina(n1618), .dinb(n718), .dout(n1619));
  jand g0978(.dina(n1619), .dinb(n1572), .dout(n1620));
  jor  g0979(.dina(n1620), .dinb(n713), .dout(n1621));
  jand g0980(.dina(n1621), .dinb(n1571), .dout(n1622));
  jor  g0981(.dina(n1622), .dinb(n708), .dout(n1623));
  jand g0982(.dina(n1623), .dinb(n1570), .dout(n1624));
  jor  g0983(.dina(n1624), .dinb(n703), .dout(n1625));
  jand g0984(.dina(n1625), .dinb(n1569), .dout(n1626));
  jor  g0985(.dina(n1626), .dinb(n698), .dout(n1627));
  jand g0986(.dina(n1627), .dinb(n1568), .dout(n1628));
  jor  g0987(.dina(n1628), .dinb(n693), .dout(n1629));
  jand g0988(.dina(n1629), .dinb(n1567), .dout(n1630));
  jor  g0989(.dina(n1630), .dinb(n688), .dout(n1631));
  jand g0990(.dina(n1631), .dinb(n1566), .dout(n1632));
  jor  g0991(.dina(n1632), .dinb(n683), .dout(n1633));
  jand g0992(.dina(n1633), .dinb(n1565), .dout(n1634));
  jor  g0993(.dina(n1634), .dinb(n678), .dout(n1635));
  jand g0994(.dina(n1635), .dinb(n1564), .dout(n1636));
  jor  g0995(.dina(n1636), .dinb(n673), .dout(n1637));
  jand g0996(.dina(n1637), .dinb(n1563), .dout(n1638));
  jor  g0997(.dina(n1638), .dinb(n668), .dout(n1639));
  jand g0998(.dina(n1639), .dinb(n1562), .dout(n1640));
  jor  g0999(.dina(n1640), .dinb(n663), .dout(n1641));
  jand g1000(.dina(n1641), .dinb(n1561), .dout(n1642));
  jor  g1001(.dina(n1642), .dinb(n658), .dout(n1643));
  jand g1002(.dina(n1643), .dinb(n1560), .dout(n1644));
  jor  g1003(.dina(n1644), .dinb(n653), .dout(n1645));
  jand g1004(.dina(n1645), .dinb(n1559), .dout(n1646));
  jor  g1005(.dina(n1646), .dinb(n648), .dout(n1647));
  jand g1006(.dina(n1647), .dinb(n1558), .dout(n1648));
  jor  g1007(.dina(n1648), .dinb(n643), .dout(n1649));
  jnot g1008(.din(n853), .dout(n1650));
  jand g1009(.dina(n1650), .dinb(n1649), .dout(n1651));
  jor  g1010(.dina(n880), .dinb(n1651), .dout(n1652));
  jnot g1011(.din(n915), .dout(n1653));
  jand g1012(.dina(n1653), .dinb(n1652), .dout(n1654));
  jor  g1013(.dina(n939), .dinb(n1654), .dout(n1655));
  jnot g1014(.din(n974), .dout(n1656));
  jand g1015(.dina(n1656), .dinb(n1655), .dout(n1657));
  jor  g1016(.dina(n1001), .dinb(n1657), .dout(n1658));
  jnot g1017(.din(n1032), .dout(n1659));
  jand g1018(.dina(n1659), .dinb(n1658), .dout(n1660));
  jor  g1019(.dina(n1056), .dinb(n1660), .dout(n1661));
  jnot g1020(.din(n1091), .dout(n1662));
  jand g1021(.dina(n1662), .dinb(n1661), .dout(n1663));
  jor  g1022(.dina(n1103), .dinb(n1663), .dout(n1664));
  jnot g1023(.din(n1120), .dout(n1665));
  jand g1024(.dina(n1665), .dinb(n1664), .dout(n1666));
  jor  g1025(.dina(n1132), .dinb(n1666), .dout(n1667));
  jnot g1026(.din(n1149), .dout(n1668));
  jand g1027(.dina(n1668), .dinb(n1667), .dout(n1669));
  jor  g1028(.dina(n1161), .dinb(n1669), .dout(n1670));
  jnot g1029(.din(n1178), .dout(n1671));
  jand g1030(.dina(n1671), .dinb(n1670), .dout(n1672));
  jor  g1031(.dina(n1190), .dinb(n1672), .dout(n1673));
  jnot g1032(.din(n1207), .dout(n1674));
  jand g1033(.dina(n1674), .dinb(n1673), .dout(n1675));
  jor  g1034(.dina(n1219), .dinb(n1675), .dout(n1676));
  jnot g1035(.din(n1236), .dout(n1677));
  jand g1036(.dina(n1677), .dinb(n1676), .dout(n1678));
  jor  g1037(.dina(n1248), .dinb(n1678), .dout(n1679));
  jnot g1038(.din(n1265), .dout(n1680));
  jand g1039(.dina(n1680), .dinb(n1679), .dout(n1681));
  jor  g1040(.dina(n1277), .dinb(n1681), .dout(n1682));
  jnot g1041(.din(n1294), .dout(n1683));
  jand g1042(.dina(n1683), .dinb(n1682), .dout(n1684));
  jor  g1043(.dina(n1306), .dinb(n1684), .dout(n1685));
  jnot g1044(.din(n1323), .dout(n1686));
  jand g1045(.dina(n1686), .dinb(n1685), .dout(n1687));
  jor  g1046(.dina(n1335), .dinb(n1687), .dout(n1688));
  jnot g1047(.din(n1352), .dout(n1689));
  jand g1048(.dina(n1689), .dinb(n1688), .dout(n1690));
  jor  g1049(.dina(n1364), .dinb(n1690), .dout(n1691));
  jnot g1050(.din(n1381), .dout(n1692));
  jand g1051(.dina(n1692), .dinb(n1691), .dout(n1693));
  jor  g1052(.dina(n1393), .dinb(n1693), .dout(n1694));
  jnot g1053(.din(n1410), .dout(n1695));
  jand g1054(.dina(n1695), .dinb(n1694), .dout(n1696));
  jor  g1055(.dina(n1422), .dinb(n1696), .dout(n1697));
  jnot g1056(.din(n1439), .dout(n1698));
  jand g1057(.dina(n1698), .dinb(n1697), .dout(n1699));
  jor  g1058(.dina(n1451), .dinb(n1699), .dout(n1700));
  jnot g1059(.din(n1468), .dout(n1701));
  jand g1060(.dina(n1701), .dinb(n1700), .dout(n1702));
  jor  g1061(.dina(n1480), .dinb(n1702), .dout(n1703));
  jnot g1062(.din(n1497), .dout(n1704));
  jand g1063(.dina(n1704), .dinb(n1703), .dout(n1705));
  jor  g1064(.dina(n1509), .dinb(n1705), .dout(n1706));
  jnot g1065(.din(n1526), .dout(n1707));
  jand g1066(.dina(n1707), .dinb(n1706), .dout(n1708));
  jor  g1067(.dina(n1538), .dinb(n1708), .dout(n1709));
  jnot g1068(.din(n1555), .dout(n1710));
  jand g1069(.dina(n1710), .dinb(n1709), .dout(n1711));
  jand g1070(.dina(n1711), .dinb(\in3[0] ), .dout(n1712));
  jor  g1071(.dina(n1712), .dinb(n1557), .dout(n1713));
  jnot g1072(.din(\in0[30] ), .dout(n1714));
  jand g1073(.dina(\in1[30] ), .dinb(n1714), .dout(n1715));
  jnot g1074(.din(n1715), .dout(n1716));
  jnot g1075(.din(\in1[29] ), .dout(n1717));
  jand g1076(.dina(n1717), .dinb(\in0[29] ), .dout(n1718));
  jnot g1077(.din(\in0[29] ), .dout(n1719));
  jand g1078(.dina(\in1[29] ), .dinb(n1719), .dout(n1720));
  jnot g1079(.din(n1720), .dout(n1721));
  jnot g1080(.din(\in1[28] ), .dout(n1722));
  jand g1081(.dina(n1722), .dinb(\in0[28] ), .dout(n1723));
  jnot g1082(.din(\in0[28] ), .dout(n1724));
  jand g1083(.dina(\in1[28] ), .dinb(n1724), .dout(n1725));
  jnot g1084(.din(n1725), .dout(n1726));
  jnot g1085(.din(\in1[27] ), .dout(n1727));
  jand g1086(.dina(n1727), .dinb(\in0[27] ), .dout(n1728));
  jnot g1087(.din(\in0[27] ), .dout(n1729));
  jand g1088(.dina(\in1[27] ), .dinb(n1729), .dout(n1730));
  jnot g1089(.din(n1730), .dout(n1731));
  jnot g1090(.din(\in1[26] ), .dout(n1732));
  jand g1091(.dina(n1732), .dinb(\in0[26] ), .dout(n1733));
  jnot g1092(.din(\in0[26] ), .dout(n1734));
  jand g1093(.dina(\in1[26] ), .dinb(n1734), .dout(n1735));
  jnot g1094(.din(n1735), .dout(n1736));
  jnot g1095(.din(\in1[25] ), .dout(n1737));
  jand g1096(.dina(n1737), .dinb(\in0[25] ), .dout(n1738));
  jnot g1097(.din(\in0[25] ), .dout(n1739));
  jand g1098(.dina(\in1[25] ), .dinb(n1739), .dout(n1740));
  jnot g1099(.din(n1740), .dout(n1741));
  jnot g1100(.din(\in1[24] ), .dout(n1742));
  jand g1101(.dina(n1742), .dinb(\in0[24] ), .dout(n1743));
  jnot g1102(.din(\in0[24] ), .dout(n1744));
  jand g1103(.dina(\in1[24] ), .dinb(n1744), .dout(n1745));
  jnot g1104(.din(n1745), .dout(n1746));
  jnot g1105(.din(\in1[23] ), .dout(n1747));
  jand g1106(.dina(n1747), .dinb(\in0[23] ), .dout(n1748));
  jnot g1107(.din(\in0[23] ), .dout(n1749));
  jand g1108(.dina(\in1[23] ), .dinb(n1749), .dout(n1750));
  jnot g1109(.din(n1750), .dout(n1751));
  jnot g1110(.din(\in1[22] ), .dout(n1752));
  jand g1111(.dina(n1752), .dinb(\in0[22] ), .dout(n1753));
  jnot g1112(.din(\in0[22] ), .dout(n1754));
  jand g1113(.dina(\in1[22] ), .dinb(n1754), .dout(n1755));
  jnot g1114(.din(n1755), .dout(n1756));
  jnot g1115(.din(\in1[21] ), .dout(n1757));
  jand g1116(.dina(n1757), .dinb(\in0[21] ), .dout(n1758));
  jnot g1117(.din(\in0[21] ), .dout(n1759));
  jand g1118(.dina(\in1[21] ), .dinb(n1759), .dout(n1760));
  jnot g1119(.din(n1760), .dout(n1761));
  jnot g1120(.din(\in1[20] ), .dout(n1762));
  jand g1121(.dina(n1762), .dinb(\in0[20] ), .dout(n1763));
  jnot g1122(.din(\in0[20] ), .dout(n1764));
  jand g1123(.dina(\in1[20] ), .dinb(n1764), .dout(n1765));
  jnot g1124(.din(n1765), .dout(n1766));
  jnot g1125(.din(\in1[19] ), .dout(n1767));
  jand g1126(.dina(n1767), .dinb(\in0[19] ), .dout(n1768));
  jnot g1127(.din(\in0[19] ), .dout(n1769));
  jand g1128(.dina(\in1[19] ), .dinb(n1769), .dout(n1770));
  jnot g1129(.din(n1770), .dout(n1771));
  jnot g1130(.din(\in1[18] ), .dout(n1772));
  jand g1131(.dina(n1772), .dinb(\in0[18] ), .dout(n1773));
  jnot g1132(.din(\in0[18] ), .dout(n1774));
  jand g1133(.dina(\in1[18] ), .dinb(n1774), .dout(n1775));
  jnot g1134(.din(n1775), .dout(n1776));
  jnot g1135(.din(\in1[17] ), .dout(n1777));
  jand g1136(.dina(n1777), .dinb(\in0[17] ), .dout(n1778));
  jnot g1137(.din(\in0[17] ), .dout(n1779));
  jand g1138(.dina(\in1[17] ), .dinb(n1779), .dout(n1780));
  jnot g1139(.din(n1780), .dout(n1781));
  jnot g1140(.din(\in1[16] ), .dout(n1782));
  jand g1141(.dina(n1782), .dinb(\in0[16] ), .dout(n1783));
  jnot g1142(.din(\in0[16] ), .dout(n1784));
  jand g1143(.dina(\in1[16] ), .dinb(n1784), .dout(n1785));
  jnot g1144(.din(n1785), .dout(n1786));
  jnot g1145(.din(\in1[15] ), .dout(n1787));
  jand g1146(.dina(n1787), .dinb(\in0[15] ), .dout(n1788));
  jnot g1147(.din(\in0[15] ), .dout(n1789));
  jand g1148(.dina(\in1[15] ), .dinb(n1789), .dout(n1790));
  jnot g1149(.din(n1790), .dout(n1791));
  jnot g1150(.din(\in1[14] ), .dout(n1792));
  jand g1151(.dina(n1792), .dinb(\in0[14] ), .dout(n1793));
  jnot g1152(.din(\in0[14] ), .dout(n1794));
  jand g1153(.dina(\in1[14] ), .dinb(n1794), .dout(n1795));
  jnot g1154(.din(n1795), .dout(n1796));
  jnot g1155(.din(\in1[13] ), .dout(n1797));
  jand g1156(.dina(n1797), .dinb(\in0[13] ), .dout(n1798));
  jnot g1157(.din(\in0[13] ), .dout(n1799));
  jand g1158(.dina(\in1[13] ), .dinb(n1799), .dout(n1800));
  jnot g1159(.din(n1800), .dout(n1801));
  jnot g1160(.din(\in1[12] ), .dout(n1802));
  jand g1161(.dina(n1802), .dinb(\in0[12] ), .dout(n1803));
  jnot g1162(.din(\in0[12] ), .dout(n1804));
  jand g1163(.dina(\in1[12] ), .dinb(n1804), .dout(n1805));
  jnot g1164(.din(n1805), .dout(n1806));
  jnot g1165(.din(\in1[11] ), .dout(n1807));
  jand g1166(.dina(n1807), .dinb(\in0[11] ), .dout(n1808));
  jnot g1167(.din(\in0[11] ), .dout(n1809));
  jand g1168(.dina(\in1[11] ), .dinb(n1809), .dout(n1810));
  jnot g1169(.din(n1810), .dout(n1811));
  jnot g1170(.din(\in1[10] ), .dout(n1812));
  jand g1171(.dina(n1812), .dinb(\in0[10] ), .dout(n1813));
  jnot g1172(.din(\in0[10] ), .dout(n1814));
  jand g1173(.dina(\in1[10] ), .dinb(n1814), .dout(n1815));
  jnot g1174(.din(n1815), .dout(n1816));
  jnot g1175(.din(\in1[9] ), .dout(n1817));
  jand g1176(.dina(n1817), .dinb(\in0[9] ), .dout(n1818));
  jnot g1177(.din(\in0[9] ), .dout(n1819));
  jand g1178(.dina(\in1[9] ), .dinb(n1819), .dout(n1820));
  jnot g1179(.din(n1820), .dout(n1821));
  jnot g1180(.din(\in1[8] ), .dout(n1822));
  jand g1181(.dina(n1822), .dinb(\in0[8] ), .dout(n1823));
  jnot g1182(.din(\in0[8] ), .dout(n1824));
  jand g1183(.dina(\in1[8] ), .dinb(n1824), .dout(n1825));
  jnot g1184(.din(n1825), .dout(n1826));
  jnot g1185(.din(\in1[7] ), .dout(n1827));
  jand g1186(.dina(n1827), .dinb(\in0[7] ), .dout(n1828));
  jnot g1187(.din(\in0[7] ), .dout(n1829));
  jand g1188(.dina(\in1[7] ), .dinb(n1829), .dout(n1830));
  jnot g1189(.din(n1830), .dout(n1831));
  jnot g1190(.din(\in1[6] ), .dout(n1832));
  jand g1191(.dina(n1832), .dinb(\in0[6] ), .dout(n1833));
  jnot g1192(.din(\in0[6] ), .dout(n1834));
  jand g1193(.dina(\in1[6] ), .dinb(n1834), .dout(n1835));
  jnot g1194(.din(n1835), .dout(n1836));
  jnot g1195(.din(\in1[5] ), .dout(n1837));
  jand g1196(.dina(n1837), .dinb(\in0[5] ), .dout(n1838));
  jnot g1197(.din(\in0[5] ), .dout(n1839));
  jand g1198(.dina(\in1[5] ), .dinb(n1839), .dout(n1840));
  jnot g1199(.din(n1840), .dout(n1841));
  jnot g1200(.din(\in1[4] ), .dout(n1842));
  jand g1201(.dina(n1842), .dinb(\in0[4] ), .dout(n1843));
  jnot g1202(.din(\in0[4] ), .dout(n1844));
  jand g1203(.dina(\in1[4] ), .dinb(n1844), .dout(n1845));
  jnot g1204(.din(n1845), .dout(n1846));
  jnot g1205(.din(\in1[3] ), .dout(n1847));
  jand g1206(.dina(n1847), .dinb(\in0[3] ), .dout(n1848));
  jnot g1207(.din(\in0[3] ), .dout(n1849));
  jand g1208(.dina(\in1[3] ), .dinb(n1849), .dout(n1850));
  jnot g1209(.din(n1850), .dout(n1851));
  jnot g1210(.din(\in1[2] ), .dout(n1852));
  jand g1211(.dina(n1852), .dinb(\in0[2] ), .dout(n1853));
  jnot g1212(.din(\in0[2] ), .dout(n1854));
  jand g1213(.dina(\in1[2] ), .dinb(n1854), .dout(n1855));
  jnot g1214(.din(n1855), .dout(n1856));
  jnot g1215(.din(\in1[1] ), .dout(n1857));
  jand g1216(.dina(n1857), .dinb(\in0[1] ), .dout(n1858));
  jor  g1217(.dina(n1857), .dinb(\in0[1] ), .dout(n1859));
  jnot g1218(.din(\in1[0] ), .dout(n1860));
  jand g1219(.dina(n1860), .dinb(\in0[0] ), .dout(n1861));
  jand g1220(.dina(n1861), .dinb(n1859), .dout(n1862));
  jor  g1221(.dina(n1862), .dinb(n1858), .dout(n1863));
  jand g1222(.dina(n1863), .dinb(n1856), .dout(n1864));
  jor  g1223(.dina(n1864), .dinb(n1853), .dout(n1865));
  jand g1224(.dina(n1865), .dinb(n1851), .dout(n1866));
  jor  g1225(.dina(n1866), .dinb(n1848), .dout(n1867));
  jand g1226(.dina(n1867), .dinb(n1846), .dout(n1868));
  jor  g1227(.dina(n1868), .dinb(n1843), .dout(n1869));
  jand g1228(.dina(n1869), .dinb(n1841), .dout(n1870));
  jor  g1229(.dina(n1870), .dinb(n1838), .dout(n1871));
  jand g1230(.dina(n1871), .dinb(n1836), .dout(n1872));
  jor  g1231(.dina(n1872), .dinb(n1833), .dout(n1873));
  jand g1232(.dina(n1873), .dinb(n1831), .dout(n1874));
  jor  g1233(.dina(n1874), .dinb(n1828), .dout(n1875));
  jand g1234(.dina(n1875), .dinb(n1826), .dout(n1876));
  jor  g1235(.dina(n1876), .dinb(n1823), .dout(n1877));
  jand g1236(.dina(n1877), .dinb(n1821), .dout(n1878));
  jor  g1237(.dina(n1878), .dinb(n1818), .dout(n1879));
  jand g1238(.dina(n1879), .dinb(n1816), .dout(n1880));
  jor  g1239(.dina(n1880), .dinb(n1813), .dout(n1881));
  jand g1240(.dina(n1881), .dinb(n1811), .dout(n1882));
  jor  g1241(.dina(n1882), .dinb(n1808), .dout(n1883));
  jand g1242(.dina(n1883), .dinb(n1806), .dout(n1884));
  jor  g1243(.dina(n1884), .dinb(n1803), .dout(n1885));
  jand g1244(.dina(n1885), .dinb(n1801), .dout(n1886));
  jor  g1245(.dina(n1886), .dinb(n1798), .dout(n1887));
  jand g1246(.dina(n1887), .dinb(n1796), .dout(n1888));
  jor  g1247(.dina(n1888), .dinb(n1793), .dout(n1889));
  jand g1248(.dina(n1889), .dinb(n1791), .dout(n1890));
  jor  g1249(.dina(n1890), .dinb(n1788), .dout(n1891));
  jand g1250(.dina(n1891), .dinb(n1786), .dout(n1892));
  jor  g1251(.dina(n1892), .dinb(n1783), .dout(n1893));
  jand g1252(.dina(n1893), .dinb(n1781), .dout(n1894));
  jor  g1253(.dina(n1894), .dinb(n1778), .dout(n1895));
  jand g1254(.dina(n1895), .dinb(n1776), .dout(n1896));
  jor  g1255(.dina(n1896), .dinb(n1773), .dout(n1897));
  jand g1256(.dina(n1897), .dinb(n1771), .dout(n1898));
  jor  g1257(.dina(n1898), .dinb(n1768), .dout(n1899));
  jand g1258(.dina(n1899), .dinb(n1766), .dout(n1900));
  jor  g1259(.dina(n1900), .dinb(n1763), .dout(n1901));
  jand g1260(.dina(n1901), .dinb(n1761), .dout(n1902));
  jor  g1261(.dina(n1902), .dinb(n1758), .dout(n1903));
  jand g1262(.dina(n1903), .dinb(n1756), .dout(n1904));
  jor  g1263(.dina(n1904), .dinb(n1753), .dout(n1905));
  jand g1264(.dina(n1905), .dinb(n1751), .dout(n1906));
  jor  g1265(.dina(n1906), .dinb(n1748), .dout(n1907));
  jand g1266(.dina(n1907), .dinb(n1746), .dout(n1908));
  jor  g1267(.dina(n1908), .dinb(n1743), .dout(n1909));
  jand g1268(.dina(n1909), .dinb(n1741), .dout(n1910));
  jor  g1269(.dina(n1910), .dinb(n1738), .dout(n1911));
  jand g1270(.dina(n1911), .dinb(n1736), .dout(n1912));
  jor  g1271(.dina(n1912), .dinb(n1733), .dout(n1913));
  jand g1272(.dina(n1913), .dinb(n1731), .dout(n1914));
  jor  g1273(.dina(n1914), .dinb(n1728), .dout(n1915));
  jand g1274(.dina(n1915), .dinb(n1726), .dout(n1916));
  jor  g1275(.dina(n1916), .dinb(n1723), .dout(n1917));
  jand g1276(.dina(n1917), .dinb(n1721), .dout(n1918));
  jor  g1277(.dina(n1918), .dinb(n1718), .dout(n1919));
  jand g1278(.dina(n1919), .dinb(n1716), .dout(n1920));
  jnot g1279(.din(\in1[30] ), .dout(n1921));
  jand g1280(.dina(n1921), .dinb(\in0[30] ), .dout(n1922));
  jnot g1281(.din(\in1[31] ), .dout(n1923));
  jand g1282(.dina(n1923), .dinb(\in0[31] ), .dout(n1924));
  jor  g1283(.dina(n1924), .dinb(n1922), .dout(n1925));
  jor  g1284(.dina(n1925), .dinb(n1920), .dout(n1926));
  jnot g1285(.din(\in0[37] ), .dout(n1927));
  jand g1286(.dina(\in1[37] ), .dinb(n1927), .dout(n1928));
  jnot g1287(.din(\in0[39] ), .dout(n1929));
  jand g1288(.dina(\in1[39] ), .dinb(n1929), .dout(n1930));
  jnot g1289(.din(\in0[38] ), .dout(n1931));
  jand g1290(.dina(\in1[38] ), .dinb(n1931), .dout(n1932));
  jor  g1291(.dina(n1932), .dinb(n1930), .dout(n1933));
  jor  g1292(.dina(n1933), .dinb(n1928), .dout(n1934));
  jnot g1293(.din(\in0[35] ), .dout(n1935));
  jand g1294(.dina(\in1[35] ), .dinb(n1935), .dout(n1936));
  jnot g1295(.din(\in0[34] ), .dout(n1937));
  jand g1296(.dina(\in1[34] ), .dinb(n1937), .dout(n1938));
  jor  g1297(.dina(n1938), .dinb(n1936), .dout(n1939));
  jnot g1298(.din(\in0[32] ), .dout(n1940));
  jand g1299(.dina(\in1[32] ), .dinb(n1940), .dout(n1941));
  jnot g1300(.din(\in0[33] ), .dout(n1942));
  jand g1301(.dina(\in1[33] ), .dinb(n1942), .dout(n1943));
  jor  g1302(.dina(n1943), .dinb(n1941), .dout(n1944));
  jnot g1303(.din(\in0[36] ), .dout(n1945));
  jand g1304(.dina(\in1[36] ), .dinb(n1945), .dout(n1946));
  jnot g1305(.din(\in0[31] ), .dout(n1947));
  jand g1306(.dina(\in1[31] ), .dinb(n1947), .dout(n1948));
  jor  g1307(.dina(n1948), .dinb(n1946), .dout(n1949));
  jor  g1308(.dina(n1949), .dinb(n1944), .dout(n1950));
  jor  g1309(.dina(n1950), .dinb(n1939), .dout(n1951));
  jor  g1310(.dina(n1951), .dinb(n1934), .dout(n1952));
  jnot g1311(.din(n1952), .dout(n1953));
  jand g1312(.dina(n1953), .dinb(n1926), .dout(n1954));
  jnot g1313(.din(n1934), .dout(n1955));
  jnot g1314(.din(n1946), .dout(n1956));
  jnot g1315(.din(\in1[35] ), .dout(n1957));
  jand g1316(.dina(n1957), .dinb(\in0[35] ), .dout(n1958));
  jnot g1317(.din(n1939), .dout(n1959));
  jnot g1318(.din(n1943), .dout(n1960));
  jnot g1319(.din(\in1[32] ), .dout(n1961));
  jand g1320(.dina(n1961), .dinb(\in0[32] ), .dout(n1962));
  jand g1321(.dina(n1962), .dinb(n1960), .dout(n1963));
  jnot g1322(.din(\in1[33] ), .dout(n1964));
  jand g1323(.dina(n1964), .dinb(\in0[33] ), .dout(n1965));
  jnot g1324(.din(\in1[34] ), .dout(n1966));
  jand g1325(.dina(n1966), .dinb(\in0[34] ), .dout(n1967));
  jor  g1326(.dina(n1967), .dinb(n1965), .dout(n1968));
  jor  g1327(.dina(n1968), .dinb(n1963), .dout(n1969));
  jand g1328(.dina(n1969), .dinb(n1959), .dout(n1970));
  jor  g1329(.dina(n1970), .dinb(n1958), .dout(n1971));
  jand g1330(.dina(n1971), .dinb(n1956), .dout(n1972));
  jnot g1331(.din(\in1[36] ), .dout(n1973));
  jand g1332(.dina(n1973), .dinb(\in0[36] ), .dout(n1974));
  jnot g1333(.din(\in1[37] ), .dout(n1975));
  jand g1334(.dina(n1975), .dinb(\in0[37] ), .dout(n1976));
  jor  g1335(.dina(n1976), .dinb(n1974), .dout(n1977));
  jor  g1336(.dina(n1977), .dinb(n1972), .dout(n1978));
  jand g1337(.dina(n1978), .dinb(n1955), .dout(n1979));
  jnot g1338(.din(n1930), .dout(n1980));
  jnot g1339(.din(\in1[38] ), .dout(n1981));
  jand g1340(.dina(n1981), .dinb(\in0[38] ), .dout(n1982));
  jand g1341(.dina(n1982), .dinb(n1980), .dout(n1983));
  jnot g1342(.din(\in1[39] ), .dout(n1984));
  jand g1343(.dina(n1984), .dinb(\in0[39] ), .dout(n1985));
  jor  g1344(.dina(n1985), .dinb(n1983), .dout(n1986));
  jor  g1345(.dina(n1986), .dinb(n1979), .dout(n1987));
  jor  g1346(.dina(n1987), .dinb(n1954), .dout(n1988));
  jnot g1347(.din(\in0[45] ), .dout(n1989));
  jand g1348(.dina(\in1[45] ), .dinb(n1989), .dout(n1990));
  jnot g1349(.din(\in0[47] ), .dout(n1991));
  jand g1350(.dina(\in1[47] ), .dinb(n1991), .dout(n1992));
  jnot g1351(.din(\in0[46] ), .dout(n1993));
  jand g1352(.dina(\in1[46] ), .dinb(n1993), .dout(n1994));
  jor  g1353(.dina(n1994), .dinb(n1992), .dout(n1995));
  jor  g1354(.dina(n1995), .dinb(n1990), .dout(n1996));
  jnot g1355(.din(\in0[43] ), .dout(n1997));
  jand g1356(.dina(\in1[43] ), .dinb(n1997), .dout(n1998));
  jnot g1357(.din(\in0[42] ), .dout(n1999));
  jand g1358(.dina(\in1[42] ), .dinb(n1999), .dout(n2000));
  jor  g1359(.dina(n2000), .dinb(n1998), .dout(n2001));
  jnot g1360(.din(\in0[44] ), .dout(n2002));
  jand g1361(.dina(\in1[44] ), .dinb(n2002), .dout(n2003));
  jnot g1362(.din(\in0[40] ), .dout(n2004));
  jand g1363(.dina(\in1[40] ), .dinb(n2004), .dout(n2005));
  jnot g1364(.din(\in0[41] ), .dout(n2006));
  jand g1365(.dina(\in1[41] ), .dinb(n2006), .dout(n2007));
  jor  g1366(.dina(n2007), .dinb(n2005), .dout(n2008));
  jor  g1367(.dina(n2008), .dinb(n2003), .dout(n2009));
  jor  g1368(.dina(n2009), .dinb(n2001), .dout(n2010));
  jor  g1369(.dina(n2010), .dinb(n1996), .dout(n2011));
  jnot g1370(.din(n2011), .dout(n2012));
  jand g1371(.dina(n2012), .dinb(n1988), .dout(n2013));
  jnot g1372(.din(n1996), .dout(n2014));
  jnot g1373(.din(n2003), .dout(n2015));
  jnot g1374(.din(\in1[43] ), .dout(n2016));
  jand g1375(.dina(n2016), .dinb(\in0[43] ), .dout(n2017));
  jnot g1376(.din(n2001), .dout(n2018));
  jnot g1377(.din(n2007), .dout(n2019));
  jnot g1378(.din(\in1[40] ), .dout(n2020));
  jand g1379(.dina(n2020), .dinb(\in0[40] ), .dout(n2021));
  jand g1380(.dina(n2021), .dinb(n2019), .dout(n2022));
  jnot g1381(.din(\in1[41] ), .dout(n2023));
  jand g1382(.dina(n2023), .dinb(\in0[41] ), .dout(n2024));
  jnot g1383(.din(\in1[42] ), .dout(n2025));
  jand g1384(.dina(n2025), .dinb(\in0[42] ), .dout(n2026));
  jor  g1385(.dina(n2026), .dinb(n2024), .dout(n2027));
  jor  g1386(.dina(n2027), .dinb(n2022), .dout(n2028));
  jand g1387(.dina(n2028), .dinb(n2018), .dout(n2029));
  jor  g1388(.dina(n2029), .dinb(n2017), .dout(n2030));
  jand g1389(.dina(n2030), .dinb(n2015), .dout(n2031));
  jnot g1390(.din(\in1[44] ), .dout(n2032));
  jand g1391(.dina(n2032), .dinb(\in0[44] ), .dout(n2033));
  jnot g1392(.din(\in1[45] ), .dout(n2034));
  jand g1393(.dina(n2034), .dinb(\in0[45] ), .dout(n2035));
  jor  g1394(.dina(n2035), .dinb(n2033), .dout(n2036));
  jor  g1395(.dina(n2036), .dinb(n2031), .dout(n2037));
  jand g1396(.dina(n2037), .dinb(n2014), .dout(n2038));
  jnot g1397(.din(n1992), .dout(n2039));
  jnot g1398(.din(\in1[46] ), .dout(n2040));
  jand g1399(.dina(n2040), .dinb(\in0[46] ), .dout(n2041));
  jand g1400(.dina(n2041), .dinb(n2039), .dout(n2042));
  jnot g1401(.din(\in1[47] ), .dout(n2043));
  jand g1402(.dina(n2043), .dinb(\in0[47] ), .dout(n2044));
  jor  g1403(.dina(n2044), .dinb(n2042), .dout(n2045));
  jor  g1404(.dina(n2045), .dinb(n2038), .dout(n2046));
  jor  g1405(.dina(n2046), .dinb(n2013), .dout(n2047));
  jnot g1406(.din(\in1[52] ), .dout(n2048));
  jnot g1407(.din(\in0[53] ), .dout(n2049));
  jand g1408(.dina(\in1[53] ), .dinb(n2049), .dout(n2050));
  jnot g1409(.din(n2050), .dout(n2051));
  jand g1410(.dina(n2051), .dinb(n2048), .dout(n2052));
  jand g1411(.dina(n2051), .dinb(\in0[52] ), .dout(n2053));
  jor  g1412(.dina(n2053), .dinb(n2052), .dout(n2054));
  jnot g1413(.din(n2054), .dout(n2055));
  jnot g1414(.din(\in0[55] ), .dout(n2056));
  jand g1415(.dina(\in1[55] ), .dinb(n2056), .dout(n2057));
  jnot g1416(.din(\in0[54] ), .dout(n2058));
  jand g1417(.dina(\in1[54] ), .dinb(n2058), .dout(n2059));
  jor  g1418(.dina(n2059), .dinb(n2057), .dout(n2060));
  jnot g1419(.din(\in0[51] ), .dout(n2061));
  jand g1420(.dina(\in1[51] ), .dinb(n2061), .dout(n2062));
  jnot g1421(.din(\in0[50] ), .dout(n2063));
  jand g1422(.dina(\in1[50] ), .dinb(n2063), .dout(n2064));
  jor  g1423(.dina(n2064), .dinb(n2062), .dout(n2065));
  jnot g1424(.din(\in0[48] ), .dout(n2066));
  jand g1425(.dina(\in1[48] ), .dinb(n2066), .dout(n2067));
  jnot g1426(.din(\in0[49] ), .dout(n2068));
  jand g1427(.dina(\in1[49] ), .dinb(n2068), .dout(n2069));
  jor  g1428(.dina(n2069), .dinb(n2067), .dout(n2070));
  jor  g1429(.dina(n2070), .dinb(n2065), .dout(n2071));
  jor  g1430(.dina(n2071), .dinb(n2060), .dout(n2072));
  jor  g1431(.dina(n2072), .dinb(n2055), .dout(n2073));
  jnot g1432(.din(n2073), .dout(n2074));
  jand g1433(.dina(n2074), .dinb(n2047), .dout(n2075));
  jnot g1434(.din(\in1[55] ), .dout(n2076));
  jand g1435(.dina(n2076), .dinb(\in0[55] ), .dout(n2077));
  jnot g1436(.din(n2060), .dout(n2078));
  jnot g1437(.din(\in1[51] ), .dout(n2079));
  jand g1438(.dina(n2079), .dinb(\in0[51] ), .dout(n2080));
  jnot g1439(.din(n2065), .dout(n2081));
  jnot g1440(.din(n2069), .dout(n2082));
  jnot g1441(.din(\in1[48] ), .dout(n2083));
  jand g1442(.dina(n2083), .dinb(\in0[48] ), .dout(n2084));
  jand g1443(.dina(n2084), .dinb(n2082), .dout(n2085));
  jnot g1444(.din(\in1[49] ), .dout(n2086));
  jand g1445(.dina(n2086), .dinb(\in0[49] ), .dout(n2087));
  jnot g1446(.din(\in1[50] ), .dout(n2088));
  jand g1447(.dina(n2088), .dinb(\in0[50] ), .dout(n2089));
  jor  g1448(.dina(n2089), .dinb(n2087), .dout(n2090));
  jor  g1449(.dina(n2090), .dinb(n2085), .dout(n2091));
  jand g1450(.dina(n2091), .dinb(n2081), .dout(n2092));
  jor  g1451(.dina(n2092), .dinb(n2080), .dout(n2093));
  jand g1452(.dina(n2093), .dinb(n2054), .dout(n2094));
  jand g1453(.dina(n2052), .dinb(\in0[52] ), .dout(n2095));
  jnot g1454(.din(\in1[53] ), .dout(n2096));
  jand g1455(.dina(n2096), .dinb(\in0[53] ), .dout(n2097));
  jnot g1456(.din(\in1[54] ), .dout(n2098));
  jand g1457(.dina(n2098), .dinb(\in0[54] ), .dout(n2099));
  jor  g1458(.dina(n2099), .dinb(n2097), .dout(n2100));
  jor  g1459(.dina(n2100), .dinb(n2095), .dout(n2101));
  jor  g1460(.dina(n2101), .dinb(n2094), .dout(n2102));
  jand g1461(.dina(n2102), .dinb(n2078), .dout(n2103));
  jor  g1462(.dina(n2103), .dinb(n2077), .dout(n2104));
  jor  g1463(.dina(n2104), .dinb(n2075), .dout(n2105));
  jnot g1464(.din(\in0[61] ), .dout(n2106));
  jand g1465(.dina(\in1[61] ), .dinb(n2106), .dout(n2107));
  jnot g1466(.din(\in0[63] ), .dout(n2108));
  jand g1467(.dina(\in1[63] ), .dinb(n2108), .dout(n2109));
  jnot g1468(.din(\in0[62] ), .dout(n2110));
  jand g1469(.dina(\in1[62] ), .dinb(n2110), .dout(n2111));
  jor  g1470(.dina(n2111), .dinb(n2109), .dout(n2112));
  jor  g1471(.dina(n2112), .dinb(n2107), .dout(n2113));
  jnot g1472(.din(\in0[59] ), .dout(n2114));
  jand g1473(.dina(\in1[59] ), .dinb(n2114), .dout(n2115));
  jnot g1474(.din(\in0[58] ), .dout(n2116));
  jand g1475(.dina(\in1[58] ), .dinb(n2116), .dout(n2117));
  jor  g1476(.dina(n2117), .dinb(n2115), .dout(n2118));
  jnot g1477(.din(\in0[60] ), .dout(n2119));
  jand g1478(.dina(\in1[60] ), .dinb(n2119), .dout(n2120));
  jnot g1479(.din(\in0[56] ), .dout(n2121));
  jand g1480(.dina(\in1[56] ), .dinb(n2121), .dout(n2122));
  jnot g1481(.din(\in0[57] ), .dout(n2123));
  jand g1482(.dina(\in1[57] ), .dinb(n2123), .dout(n2124));
  jor  g1483(.dina(n2124), .dinb(n2122), .dout(n2125));
  jor  g1484(.dina(n2125), .dinb(n2120), .dout(n2126));
  jor  g1485(.dina(n2126), .dinb(n2118), .dout(n2127));
  jor  g1486(.dina(n2127), .dinb(n2113), .dout(n2128));
  jnot g1487(.din(n2128), .dout(n2129));
  jand g1488(.dina(n2129), .dinb(n2105), .dout(n2130));
  jnot g1489(.din(n2113), .dout(n2131));
  jnot g1490(.din(n2120), .dout(n2132));
  jnot g1491(.din(\in1[59] ), .dout(n2133));
  jand g1492(.dina(n2133), .dinb(\in0[59] ), .dout(n2134));
  jnot g1493(.din(n2118), .dout(n2135));
  jnot g1494(.din(n2124), .dout(n2136));
  jnot g1495(.din(\in1[56] ), .dout(n2137));
  jand g1496(.dina(n2137), .dinb(\in0[56] ), .dout(n2138));
  jand g1497(.dina(n2138), .dinb(n2136), .dout(n2139));
  jnot g1498(.din(\in1[57] ), .dout(n2140));
  jand g1499(.dina(n2140), .dinb(\in0[57] ), .dout(n2141));
  jnot g1500(.din(\in1[58] ), .dout(n2142));
  jand g1501(.dina(n2142), .dinb(\in0[58] ), .dout(n2143));
  jor  g1502(.dina(n2143), .dinb(n2141), .dout(n2144));
  jor  g1503(.dina(n2144), .dinb(n2139), .dout(n2145));
  jand g1504(.dina(n2145), .dinb(n2135), .dout(n2146));
  jor  g1505(.dina(n2146), .dinb(n2134), .dout(n2147));
  jand g1506(.dina(n2147), .dinb(n2132), .dout(n2148));
  jnot g1507(.din(\in1[60] ), .dout(n2149));
  jand g1508(.dina(n2149), .dinb(\in0[60] ), .dout(n2150));
  jnot g1509(.din(\in1[61] ), .dout(n2151));
  jand g1510(.dina(n2151), .dinb(\in0[61] ), .dout(n2152));
  jor  g1511(.dina(n2152), .dinb(n2150), .dout(n2153));
  jor  g1512(.dina(n2153), .dinb(n2148), .dout(n2154));
  jand g1513(.dina(n2154), .dinb(n2131), .dout(n2155));
  jnot g1514(.din(n2109), .dout(n2156));
  jnot g1515(.din(\in1[62] ), .dout(n2157));
  jand g1516(.dina(n2157), .dinb(\in0[62] ), .dout(n2158));
  jand g1517(.dina(n2158), .dinb(n2156), .dout(n2159));
  jnot g1518(.din(\in1[63] ), .dout(n2160));
  jand g1519(.dina(n2160), .dinb(\in0[63] ), .dout(n2161));
  jor  g1520(.dina(n2161), .dinb(n2159), .dout(n2162));
  jor  g1521(.dina(n2162), .dinb(n2155), .dout(n2163));
  jor  g1522(.dina(n2163), .dinb(n2130), .dout(n2164));
  jnot g1523(.din(\in0[67] ), .dout(n2165));
  jand g1524(.dina(\in1[67] ), .dinb(n2165), .dout(n2166));
  jnot g1525(.din(\in0[66] ), .dout(n2167));
  jand g1526(.dina(\in1[66] ), .dinb(n2167), .dout(n2168));
  jor  g1527(.dina(n2168), .dinb(n2166), .dout(n2169));
  jnot g1528(.din(\in0[65] ), .dout(n2170));
  jand g1529(.dina(\in1[65] ), .dinb(n2170), .dout(n2171));
  jnot g1530(.din(\in0[64] ), .dout(n2172));
  jand g1531(.dina(\in1[64] ), .dinb(n2172), .dout(n2173));
  jor  g1532(.dina(n2173), .dinb(n2171), .dout(n2174));
  jor  g1533(.dina(n2174), .dinb(n2169), .dout(n2175));
  jnot g1534(.din(n2175), .dout(n2176));
  jand g1535(.dina(n2176), .dinb(n2164), .dout(n2177));
  jnot g1536(.din(\in1[67] ), .dout(n2178));
  jand g1537(.dina(n2178), .dinb(\in0[67] ), .dout(n2179));
  jnot g1538(.din(n2169), .dout(n2180));
  jnot g1539(.din(n2171), .dout(n2181));
  jnot g1540(.din(\in1[64] ), .dout(n2182));
  jand g1541(.dina(n2182), .dinb(\in0[64] ), .dout(n2183));
  jand g1542(.dina(n2183), .dinb(n2181), .dout(n2184));
  jnot g1543(.din(\in1[65] ), .dout(n2185));
  jand g1544(.dina(n2185), .dinb(\in0[65] ), .dout(n2186));
  jnot g1545(.din(\in1[66] ), .dout(n2187));
  jand g1546(.dina(n2187), .dinb(\in0[66] ), .dout(n2188));
  jor  g1547(.dina(n2188), .dinb(n2186), .dout(n2189));
  jor  g1548(.dina(n2189), .dinb(n2184), .dout(n2190));
  jand g1549(.dina(n2190), .dinb(n2180), .dout(n2191));
  jor  g1550(.dina(n2191), .dinb(n2179), .dout(n2192));
  jor  g1551(.dina(n2192), .dinb(n2177), .dout(n2193));
  jnot g1552(.din(\in0[68] ), .dout(n2194));
  jand g1553(.dina(\in1[68] ), .dinb(n2194), .dout(n2195));
  jnot g1554(.din(\in0[69] ), .dout(n2196));
  jand g1555(.dina(\in1[69] ), .dinb(n2196), .dout(n2197));
  jnot g1556(.din(\in0[71] ), .dout(n2198));
  jand g1557(.dina(\in1[71] ), .dinb(n2198), .dout(n2199));
  jnot g1558(.din(\in0[70] ), .dout(n2200));
  jand g1559(.dina(\in1[70] ), .dinb(n2200), .dout(n2201));
  jor  g1560(.dina(n2201), .dinb(n2199), .dout(n2202));
  jor  g1561(.dina(n2202), .dinb(n2197), .dout(n2203));
  jor  g1562(.dina(n2203), .dinb(n2195), .dout(n2204));
  jnot g1563(.din(n2204), .dout(n2205));
  jand g1564(.dina(n2205), .dinb(n2193), .dout(n2206));
  jnot g1565(.din(n2203), .dout(n2207));
  jnot g1566(.din(\in1[69] ), .dout(n2208));
  jand g1567(.dina(n2208), .dinb(\in0[69] ), .dout(n2209));
  jnot g1568(.din(\in1[68] ), .dout(n2210));
  jand g1569(.dina(n2210), .dinb(\in0[68] ), .dout(n2211));
  jor  g1570(.dina(n2211), .dinb(n2209), .dout(n2212));
  jand g1571(.dina(n2212), .dinb(n2207), .dout(n2213));
  jnot g1572(.din(\in1[71] ), .dout(n2214));
  jand g1573(.dina(n2214), .dinb(\in0[71] ), .dout(n2215));
  jnot g1574(.din(n2199), .dout(n2216));
  jnot g1575(.din(\in1[70] ), .dout(n2217));
  jand g1576(.dina(n2217), .dinb(\in0[70] ), .dout(n2218));
  jand g1577(.dina(n2218), .dinb(n2216), .dout(n2219));
  jor  g1578(.dina(n2219), .dinb(n2215), .dout(n2220));
  jor  g1579(.dina(n2220), .dinb(n2213), .dout(n2221));
  jor  g1580(.dina(n2221), .dinb(n2206), .dout(n2222));
  jnot g1581(.din(\in0[75] ), .dout(n2223));
  jand g1582(.dina(\in1[75] ), .dinb(n2223), .dout(n2224));
  jnot g1583(.din(\in0[74] ), .dout(n2225));
  jand g1584(.dina(\in1[74] ), .dinb(n2225), .dout(n2226));
  jor  g1585(.dina(n2226), .dinb(n2224), .dout(n2227));
  jnot g1586(.din(\in0[73] ), .dout(n2228));
  jand g1587(.dina(\in1[73] ), .dinb(n2228), .dout(n2229));
  jnot g1588(.din(\in0[72] ), .dout(n2230));
  jand g1589(.dina(\in1[72] ), .dinb(n2230), .dout(n2231));
  jor  g1590(.dina(n2231), .dinb(n2229), .dout(n2232));
  jor  g1591(.dina(n2232), .dinb(n2227), .dout(n2233));
  jnot g1592(.din(n2233), .dout(n2234));
  jand g1593(.dina(n2234), .dinb(n2222), .dout(n2235));
  jnot g1594(.din(\in1[75] ), .dout(n2236));
  jand g1595(.dina(n2236), .dinb(\in0[75] ), .dout(n2237));
  jnot g1596(.din(n2227), .dout(n2238));
  jnot g1597(.din(n2229), .dout(n2239));
  jnot g1598(.din(\in1[72] ), .dout(n2240));
  jand g1599(.dina(n2240), .dinb(\in0[72] ), .dout(n2241));
  jand g1600(.dina(n2241), .dinb(n2239), .dout(n2242));
  jnot g1601(.din(\in1[73] ), .dout(n2243));
  jand g1602(.dina(n2243), .dinb(\in0[73] ), .dout(n2244));
  jnot g1603(.din(\in1[74] ), .dout(n2245));
  jand g1604(.dina(n2245), .dinb(\in0[74] ), .dout(n2246));
  jor  g1605(.dina(n2246), .dinb(n2244), .dout(n2247));
  jor  g1606(.dina(n2247), .dinb(n2242), .dout(n2248));
  jand g1607(.dina(n2248), .dinb(n2238), .dout(n2249));
  jor  g1608(.dina(n2249), .dinb(n2237), .dout(n2250));
  jor  g1609(.dina(n2250), .dinb(n2235), .dout(n2251));
  jnot g1610(.din(\in0[76] ), .dout(n2252));
  jand g1611(.dina(\in1[76] ), .dinb(n2252), .dout(n2253));
  jnot g1612(.din(\in0[77] ), .dout(n2254));
  jand g1613(.dina(\in1[77] ), .dinb(n2254), .dout(n2255));
  jnot g1614(.din(\in0[79] ), .dout(n2256));
  jand g1615(.dina(\in1[79] ), .dinb(n2256), .dout(n2257));
  jnot g1616(.din(\in0[78] ), .dout(n2258));
  jand g1617(.dina(\in1[78] ), .dinb(n2258), .dout(n2259));
  jor  g1618(.dina(n2259), .dinb(n2257), .dout(n2260));
  jor  g1619(.dina(n2260), .dinb(n2255), .dout(n2261));
  jor  g1620(.dina(n2261), .dinb(n2253), .dout(n2262));
  jnot g1621(.din(n2262), .dout(n2263));
  jand g1622(.dina(n2263), .dinb(n2251), .dout(n2264));
  jnot g1623(.din(n2261), .dout(n2265));
  jnot g1624(.din(\in1[77] ), .dout(n2266));
  jand g1625(.dina(n2266), .dinb(\in0[77] ), .dout(n2267));
  jnot g1626(.din(\in1[76] ), .dout(n2268));
  jand g1627(.dina(n2268), .dinb(\in0[76] ), .dout(n2269));
  jor  g1628(.dina(n2269), .dinb(n2267), .dout(n2270));
  jand g1629(.dina(n2270), .dinb(n2265), .dout(n2271));
  jnot g1630(.din(\in1[79] ), .dout(n2272));
  jand g1631(.dina(n2272), .dinb(\in0[79] ), .dout(n2273));
  jnot g1632(.din(n2257), .dout(n2274));
  jnot g1633(.din(\in1[78] ), .dout(n2275));
  jand g1634(.dina(n2275), .dinb(\in0[78] ), .dout(n2276));
  jand g1635(.dina(n2276), .dinb(n2274), .dout(n2277));
  jor  g1636(.dina(n2277), .dinb(n2273), .dout(n2278));
  jor  g1637(.dina(n2278), .dinb(n2271), .dout(n2279));
  jor  g1638(.dina(n2279), .dinb(n2264), .dout(n2280));
  jnot g1639(.din(\in0[83] ), .dout(n2281));
  jand g1640(.dina(\in1[83] ), .dinb(n2281), .dout(n2282));
  jnot g1641(.din(\in0[82] ), .dout(n2283));
  jand g1642(.dina(\in1[82] ), .dinb(n2283), .dout(n2284));
  jor  g1643(.dina(n2284), .dinb(n2282), .dout(n2285));
  jnot g1644(.din(\in0[81] ), .dout(n2286));
  jand g1645(.dina(\in1[81] ), .dinb(n2286), .dout(n2287));
  jnot g1646(.din(\in0[80] ), .dout(n2288));
  jand g1647(.dina(\in1[80] ), .dinb(n2288), .dout(n2289));
  jor  g1648(.dina(n2289), .dinb(n2287), .dout(n2290));
  jor  g1649(.dina(n2290), .dinb(n2285), .dout(n2291));
  jnot g1650(.din(n2291), .dout(n2292));
  jand g1651(.dina(n2292), .dinb(n2280), .dout(n2293));
  jnot g1652(.din(\in1[83] ), .dout(n2294));
  jand g1653(.dina(n2294), .dinb(\in0[83] ), .dout(n2295));
  jnot g1654(.din(n2285), .dout(n2296));
  jnot g1655(.din(n2287), .dout(n2297));
  jnot g1656(.din(\in1[80] ), .dout(n2298));
  jand g1657(.dina(n2298), .dinb(\in0[80] ), .dout(n2299));
  jand g1658(.dina(n2299), .dinb(n2297), .dout(n2300));
  jnot g1659(.din(\in1[81] ), .dout(n2301));
  jand g1660(.dina(n2301), .dinb(\in0[81] ), .dout(n2302));
  jnot g1661(.din(\in1[82] ), .dout(n2303));
  jand g1662(.dina(n2303), .dinb(\in0[82] ), .dout(n2304));
  jor  g1663(.dina(n2304), .dinb(n2302), .dout(n2305));
  jor  g1664(.dina(n2305), .dinb(n2300), .dout(n2306));
  jand g1665(.dina(n2306), .dinb(n2296), .dout(n2307));
  jor  g1666(.dina(n2307), .dinb(n2295), .dout(n2308));
  jor  g1667(.dina(n2308), .dinb(n2293), .dout(n2309));
  jnot g1668(.din(\in0[84] ), .dout(n2310));
  jand g1669(.dina(\in1[84] ), .dinb(n2310), .dout(n2311));
  jnot g1670(.din(\in0[85] ), .dout(n2312));
  jand g1671(.dina(\in1[85] ), .dinb(n2312), .dout(n2313));
  jnot g1672(.din(\in0[87] ), .dout(n2314));
  jand g1673(.dina(\in1[87] ), .dinb(n2314), .dout(n2315));
  jnot g1674(.din(\in0[86] ), .dout(n2316));
  jand g1675(.dina(\in1[86] ), .dinb(n2316), .dout(n2317));
  jor  g1676(.dina(n2317), .dinb(n2315), .dout(n2318));
  jor  g1677(.dina(n2318), .dinb(n2313), .dout(n2319));
  jor  g1678(.dina(n2319), .dinb(n2311), .dout(n2320));
  jnot g1679(.din(n2320), .dout(n2321));
  jand g1680(.dina(n2321), .dinb(n2309), .dout(n2322));
  jnot g1681(.din(n2319), .dout(n2323));
  jnot g1682(.din(\in1[85] ), .dout(n2324));
  jand g1683(.dina(n2324), .dinb(\in0[85] ), .dout(n2325));
  jnot g1684(.din(\in1[84] ), .dout(n2326));
  jand g1685(.dina(n2326), .dinb(\in0[84] ), .dout(n2327));
  jor  g1686(.dina(n2327), .dinb(n2325), .dout(n2328));
  jand g1687(.dina(n2328), .dinb(n2323), .dout(n2329));
  jnot g1688(.din(\in1[87] ), .dout(n2330));
  jand g1689(.dina(n2330), .dinb(\in0[87] ), .dout(n2331));
  jnot g1690(.din(n2315), .dout(n2332));
  jnot g1691(.din(\in1[86] ), .dout(n2333));
  jand g1692(.dina(n2333), .dinb(\in0[86] ), .dout(n2334));
  jand g1693(.dina(n2334), .dinb(n2332), .dout(n2335));
  jor  g1694(.dina(n2335), .dinb(n2331), .dout(n2336));
  jor  g1695(.dina(n2336), .dinb(n2329), .dout(n2337));
  jor  g1696(.dina(n2337), .dinb(n2322), .dout(n2338));
  jnot g1697(.din(\in0[91] ), .dout(n2339));
  jand g1698(.dina(\in1[91] ), .dinb(n2339), .dout(n2340));
  jnot g1699(.din(\in0[90] ), .dout(n2341));
  jand g1700(.dina(\in1[90] ), .dinb(n2341), .dout(n2342));
  jor  g1701(.dina(n2342), .dinb(n2340), .dout(n2343));
  jnot g1702(.din(\in0[89] ), .dout(n2344));
  jand g1703(.dina(\in1[89] ), .dinb(n2344), .dout(n2345));
  jnot g1704(.din(\in0[88] ), .dout(n2346));
  jand g1705(.dina(\in1[88] ), .dinb(n2346), .dout(n2347));
  jor  g1706(.dina(n2347), .dinb(n2345), .dout(n2348));
  jor  g1707(.dina(n2348), .dinb(n2343), .dout(n2349));
  jnot g1708(.din(n2349), .dout(n2350));
  jand g1709(.dina(n2350), .dinb(n2338), .dout(n2351));
  jnot g1710(.din(\in1[91] ), .dout(n2352));
  jand g1711(.dina(n2352), .dinb(\in0[91] ), .dout(n2353));
  jnot g1712(.din(n2343), .dout(n2354));
  jnot g1713(.din(n2345), .dout(n2355));
  jnot g1714(.din(\in1[88] ), .dout(n2356));
  jand g1715(.dina(n2356), .dinb(\in0[88] ), .dout(n2357));
  jand g1716(.dina(n2357), .dinb(n2355), .dout(n2358));
  jnot g1717(.din(\in1[89] ), .dout(n2359));
  jand g1718(.dina(n2359), .dinb(\in0[89] ), .dout(n2360));
  jnot g1719(.din(\in1[90] ), .dout(n2361));
  jand g1720(.dina(n2361), .dinb(\in0[90] ), .dout(n2362));
  jor  g1721(.dina(n2362), .dinb(n2360), .dout(n2363));
  jor  g1722(.dina(n2363), .dinb(n2358), .dout(n2364));
  jand g1723(.dina(n2364), .dinb(n2354), .dout(n2365));
  jor  g1724(.dina(n2365), .dinb(n2353), .dout(n2366));
  jor  g1725(.dina(n2366), .dinb(n2351), .dout(n2367));
  jnot g1726(.din(\in0[92] ), .dout(n2368));
  jand g1727(.dina(\in1[92] ), .dinb(n2368), .dout(n2369));
  jnot g1728(.din(\in0[93] ), .dout(n2370));
  jand g1729(.dina(\in1[93] ), .dinb(n2370), .dout(n2371));
  jnot g1730(.din(\in0[95] ), .dout(n2372));
  jand g1731(.dina(\in1[95] ), .dinb(n2372), .dout(n2373));
  jnot g1732(.din(\in0[94] ), .dout(n2374));
  jand g1733(.dina(\in1[94] ), .dinb(n2374), .dout(n2375));
  jor  g1734(.dina(n2375), .dinb(n2373), .dout(n2376));
  jor  g1735(.dina(n2376), .dinb(n2371), .dout(n2377));
  jor  g1736(.dina(n2377), .dinb(n2369), .dout(n2378));
  jnot g1737(.din(n2378), .dout(n2379));
  jand g1738(.dina(n2379), .dinb(n2367), .dout(n2380));
  jnot g1739(.din(n2377), .dout(n2381));
  jnot g1740(.din(\in1[93] ), .dout(n2382));
  jand g1741(.dina(n2382), .dinb(\in0[93] ), .dout(n2383));
  jnot g1742(.din(\in1[92] ), .dout(n2384));
  jand g1743(.dina(n2384), .dinb(\in0[92] ), .dout(n2385));
  jor  g1744(.dina(n2385), .dinb(n2383), .dout(n2386));
  jand g1745(.dina(n2386), .dinb(n2381), .dout(n2387));
  jnot g1746(.din(\in1[95] ), .dout(n2388));
  jand g1747(.dina(n2388), .dinb(\in0[95] ), .dout(n2389));
  jnot g1748(.din(n2373), .dout(n2390));
  jnot g1749(.din(\in1[94] ), .dout(n2391));
  jand g1750(.dina(n2391), .dinb(\in0[94] ), .dout(n2392));
  jand g1751(.dina(n2392), .dinb(n2390), .dout(n2393));
  jor  g1752(.dina(n2393), .dinb(n2389), .dout(n2394));
  jor  g1753(.dina(n2394), .dinb(n2387), .dout(n2395));
  jor  g1754(.dina(n2395), .dinb(n2380), .dout(n2396));
  jnot g1755(.din(\in0[99] ), .dout(n2397));
  jand g1756(.dina(\in1[99] ), .dinb(n2397), .dout(n2398));
  jnot g1757(.din(\in0[98] ), .dout(n2399));
  jand g1758(.dina(\in1[98] ), .dinb(n2399), .dout(n2400));
  jor  g1759(.dina(n2400), .dinb(n2398), .dout(n2401));
  jnot g1760(.din(\in0[97] ), .dout(n2402));
  jand g1761(.dina(\in1[97] ), .dinb(n2402), .dout(n2403));
  jnot g1762(.din(\in0[96] ), .dout(n2404));
  jand g1763(.dina(\in1[96] ), .dinb(n2404), .dout(n2405));
  jor  g1764(.dina(n2405), .dinb(n2403), .dout(n2406));
  jor  g1765(.dina(n2406), .dinb(n2401), .dout(n2407));
  jnot g1766(.din(n2407), .dout(n2408));
  jand g1767(.dina(n2408), .dinb(n2396), .dout(n2409));
  jnot g1768(.din(\in1[99] ), .dout(n2410));
  jand g1769(.dina(n2410), .dinb(\in0[99] ), .dout(n2411));
  jnot g1770(.din(n2401), .dout(n2412));
  jnot g1771(.din(n2403), .dout(n2413));
  jnot g1772(.din(\in1[96] ), .dout(n2414));
  jand g1773(.dina(n2414), .dinb(\in0[96] ), .dout(n2415));
  jand g1774(.dina(n2415), .dinb(n2413), .dout(n2416));
  jnot g1775(.din(\in1[97] ), .dout(n2417));
  jand g1776(.dina(n2417), .dinb(\in0[97] ), .dout(n2418));
  jnot g1777(.din(\in1[98] ), .dout(n2419));
  jand g1778(.dina(n2419), .dinb(\in0[98] ), .dout(n2420));
  jor  g1779(.dina(n2420), .dinb(n2418), .dout(n2421));
  jor  g1780(.dina(n2421), .dinb(n2416), .dout(n2422));
  jand g1781(.dina(n2422), .dinb(n2412), .dout(n2423));
  jor  g1782(.dina(n2423), .dinb(n2411), .dout(n2424));
  jor  g1783(.dina(n2424), .dinb(n2409), .dout(n2425));
  jnot g1784(.din(\in0[100] ), .dout(n2426));
  jand g1785(.dina(\in1[100] ), .dinb(n2426), .dout(n2427));
  jnot g1786(.din(\in0[101] ), .dout(n2428));
  jand g1787(.dina(\in1[101] ), .dinb(n2428), .dout(n2429));
  jnot g1788(.din(\in0[103] ), .dout(n2430));
  jand g1789(.dina(\in1[103] ), .dinb(n2430), .dout(n2431));
  jnot g1790(.din(\in0[102] ), .dout(n2432));
  jand g1791(.dina(\in1[102] ), .dinb(n2432), .dout(n2433));
  jor  g1792(.dina(n2433), .dinb(n2431), .dout(n2434));
  jor  g1793(.dina(n2434), .dinb(n2429), .dout(n2435));
  jor  g1794(.dina(n2435), .dinb(n2427), .dout(n2436));
  jnot g1795(.din(n2436), .dout(n2437));
  jand g1796(.dina(n2437), .dinb(n2425), .dout(n2438));
  jnot g1797(.din(n2435), .dout(n2439));
  jnot g1798(.din(\in1[101] ), .dout(n2440));
  jand g1799(.dina(n2440), .dinb(\in0[101] ), .dout(n2441));
  jnot g1800(.din(\in1[100] ), .dout(n2442));
  jand g1801(.dina(n2442), .dinb(\in0[100] ), .dout(n2443));
  jor  g1802(.dina(n2443), .dinb(n2441), .dout(n2444));
  jand g1803(.dina(n2444), .dinb(n2439), .dout(n2445));
  jnot g1804(.din(\in1[103] ), .dout(n2446));
  jand g1805(.dina(n2446), .dinb(\in0[103] ), .dout(n2447));
  jnot g1806(.din(n2431), .dout(n2448));
  jnot g1807(.din(\in1[102] ), .dout(n2449));
  jand g1808(.dina(n2449), .dinb(\in0[102] ), .dout(n2450));
  jand g1809(.dina(n2450), .dinb(n2448), .dout(n2451));
  jor  g1810(.dina(n2451), .dinb(n2447), .dout(n2452));
  jor  g1811(.dina(n2452), .dinb(n2445), .dout(n2453));
  jor  g1812(.dina(n2453), .dinb(n2438), .dout(n2454));
  jnot g1813(.din(\in0[107] ), .dout(n2455));
  jand g1814(.dina(\in1[107] ), .dinb(n2455), .dout(n2456));
  jnot g1815(.din(\in0[106] ), .dout(n2457));
  jand g1816(.dina(\in1[106] ), .dinb(n2457), .dout(n2458));
  jor  g1817(.dina(n2458), .dinb(n2456), .dout(n2459));
  jnot g1818(.din(\in0[105] ), .dout(n2460));
  jand g1819(.dina(\in1[105] ), .dinb(n2460), .dout(n2461));
  jnot g1820(.din(\in0[104] ), .dout(n2462));
  jand g1821(.dina(\in1[104] ), .dinb(n2462), .dout(n2463));
  jor  g1822(.dina(n2463), .dinb(n2461), .dout(n2464));
  jor  g1823(.dina(n2464), .dinb(n2459), .dout(n2465));
  jnot g1824(.din(n2465), .dout(n2466));
  jand g1825(.dina(n2466), .dinb(n2454), .dout(n2467));
  jnot g1826(.din(\in1[107] ), .dout(n2468));
  jand g1827(.dina(n2468), .dinb(\in0[107] ), .dout(n2469));
  jnot g1828(.din(n2459), .dout(n2470));
  jnot g1829(.din(n2461), .dout(n2471));
  jnot g1830(.din(\in1[104] ), .dout(n2472));
  jand g1831(.dina(n2472), .dinb(\in0[104] ), .dout(n2473));
  jand g1832(.dina(n2473), .dinb(n2471), .dout(n2474));
  jnot g1833(.din(\in1[105] ), .dout(n2475));
  jand g1834(.dina(n2475), .dinb(\in0[105] ), .dout(n2476));
  jnot g1835(.din(\in1[106] ), .dout(n2477));
  jand g1836(.dina(n2477), .dinb(\in0[106] ), .dout(n2478));
  jor  g1837(.dina(n2478), .dinb(n2476), .dout(n2479));
  jor  g1838(.dina(n2479), .dinb(n2474), .dout(n2480));
  jand g1839(.dina(n2480), .dinb(n2470), .dout(n2481));
  jor  g1840(.dina(n2481), .dinb(n2469), .dout(n2482));
  jor  g1841(.dina(n2482), .dinb(n2467), .dout(n2483));
  jnot g1842(.din(\in0[108] ), .dout(n2484));
  jand g1843(.dina(\in1[108] ), .dinb(n2484), .dout(n2485));
  jnot g1844(.din(\in0[109] ), .dout(n2486));
  jand g1845(.dina(\in1[109] ), .dinb(n2486), .dout(n2487));
  jnot g1846(.din(\in0[111] ), .dout(n2488));
  jand g1847(.dina(\in1[111] ), .dinb(n2488), .dout(n2489));
  jnot g1848(.din(\in0[110] ), .dout(n2490));
  jand g1849(.dina(\in1[110] ), .dinb(n2490), .dout(n2491));
  jor  g1850(.dina(n2491), .dinb(n2489), .dout(n2492));
  jor  g1851(.dina(n2492), .dinb(n2487), .dout(n2493));
  jor  g1852(.dina(n2493), .dinb(n2485), .dout(n2494));
  jnot g1853(.din(n2494), .dout(n2495));
  jand g1854(.dina(n2495), .dinb(n2483), .dout(n2496));
  jnot g1855(.din(n2493), .dout(n2497));
  jnot g1856(.din(\in1[109] ), .dout(n2498));
  jand g1857(.dina(n2498), .dinb(\in0[109] ), .dout(n2499));
  jnot g1858(.din(\in1[108] ), .dout(n2500));
  jand g1859(.dina(n2500), .dinb(\in0[108] ), .dout(n2501));
  jor  g1860(.dina(n2501), .dinb(n2499), .dout(n2502));
  jand g1861(.dina(n2502), .dinb(n2497), .dout(n2503));
  jnot g1862(.din(\in1[111] ), .dout(n2504));
  jand g1863(.dina(n2504), .dinb(\in0[111] ), .dout(n2505));
  jnot g1864(.din(n2489), .dout(n2506));
  jnot g1865(.din(\in1[110] ), .dout(n2507));
  jand g1866(.dina(n2507), .dinb(\in0[110] ), .dout(n2508));
  jand g1867(.dina(n2508), .dinb(n2506), .dout(n2509));
  jor  g1868(.dina(n2509), .dinb(n2505), .dout(n2510));
  jor  g1869(.dina(n2510), .dinb(n2503), .dout(n2511));
  jor  g1870(.dina(n2511), .dinb(n2496), .dout(n2512));
  jnot g1871(.din(\in0[115] ), .dout(n2513));
  jand g1872(.dina(\in1[115] ), .dinb(n2513), .dout(n2514));
  jnot g1873(.din(\in0[114] ), .dout(n2515));
  jand g1874(.dina(\in1[114] ), .dinb(n2515), .dout(n2516));
  jor  g1875(.dina(n2516), .dinb(n2514), .dout(n2517));
  jnot g1876(.din(\in0[113] ), .dout(n2518));
  jand g1877(.dina(\in1[113] ), .dinb(n2518), .dout(n2519));
  jnot g1878(.din(\in0[112] ), .dout(n2520));
  jand g1879(.dina(\in1[112] ), .dinb(n2520), .dout(n2521));
  jor  g1880(.dina(n2521), .dinb(n2519), .dout(n2522));
  jor  g1881(.dina(n2522), .dinb(n2517), .dout(n2523));
  jnot g1882(.din(n2523), .dout(n2524));
  jand g1883(.dina(n2524), .dinb(n2512), .dout(n2525));
  jnot g1884(.din(\in1[115] ), .dout(n2526));
  jand g1885(.dina(n2526), .dinb(\in0[115] ), .dout(n2527));
  jnot g1886(.din(n2517), .dout(n2528));
  jnot g1887(.din(n2519), .dout(n2529));
  jnot g1888(.din(\in1[112] ), .dout(n2530));
  jand g1889(.dina(n2530), .dinb(\in0[112] ), .dout(n2531));
  jand g1890(.dina(n2531), .dinb(n2529), .dout(n2532));
  jnot g1891(.din(\in1[113] ), .dout(n2533));
  jand g1892(.dina(n2533), .dinb(\in0[113] ), .dout(n2534));
  jnot g1893(.din(\in1[114] ), .dout(n2535));
  jand g1894(.dina(n2535), .dinb(\in0[114] ), .dout(n2536));
  jor  g1895(.dina(n2536), .dinb(n2534), .dout(n2537));
  jor  g1896(.dina(n2537), .dinb(n2532), .dout(n2538));
  jand g1897(.dina(n2538), .dinb(n2528), .dout(n2539));
  jor  g1898(.dina(n2539), .dinb(n2527), .dout(n2540));
  jor  g1899(.dina(n2540), .dinb(n2525), .dout(n2541));
  jnot g1900(.din(\in0[116] ), .dout(n2542));
  jand g1901(.dina(\in1[116] ), .dinb(n2542), .dout(n2543));
  jnot g1902(.din(\in0[117] ), .dout(n2544));
  jand g1903(.dina(\in1[117] ), .dinb(n2544), .dout(n2545));
  jnot g1904(.din(\in0[119] ), .dout(n2546));
  jand g1905(.dina(\in1[119] ), .dinb(n2546), .dout(n2547));
  jnot g1906(.din(\in0[118] ), .dout(n2548));
  jand g1907(.dina(\in1[118] ), .dinb(n2548), .dout(n2549));
  jor  g1908(.dina(n2549), .dinb(n2547), .dout(n2550));
  jor  g1909(.dina(n2550), .dinb(n2545), .dout(n2551));
  jor  g1910(.dina(n2551), .dinb(n2543), .dout(n2552));
  jnot g1911(.din(n2552), .dout(n2553));
  jand g1912(.dina(n2553), .dinb(n2541), .dout(n2554));
  jnot g1913(.din(n2551), .dout(n2555));
  jnot g1914(.din(\in1[117] ), .dout(n2556));
  jand g1915(.dina(n2556), .dinb(\in0[117] ), .dout(n2557));
  jnot g1916(.din(\in1[116] ), .dout(n2558));
  jand g1917(.dina(n2558), .dinb(\in0[116] ), .dout(n2559));
  jor  g1918(.dina(n2559), .dinb(n2557), .dout(n2560));
  jand g1919(.dina(n2560), .dinb(n2555), .dout(n2561));
  jnot g1920(.din(\in1[119] ), .dout(n2562));
  jand g1921(.dina(n2562), .dinb(\in0[119] ), .dout(n2563));
  jnot g1922(.din(n2547), .dout(n2564));
  jnot g1923(.din(\in1[118] ), .dout(n2565));
  jand g1924(.dina(n2565), .dinb(\in0[118] ), .dout(n2566));
  jand g1925(.dina(n2566), .dinb(n2564), .dout(n2567));
  jor  g1926(.dina(n2567), .dinb(n2563), .dout(n2568));
  jor  g1927(.dina(n2568), .dinb(n2561), .dout(n2569));
  jor  g1928(.dina(n2569), .dinb(n2554), .dout(n2570));
  jnot g1929(.din(\in0[123] ), .dout(n2571));
  jand g1930(.dina(\in1[123] ), .dinb(n2571), .dout(n2572));
  jnot g1931(.din(\in0[122] ), .dout(n2573));
  jand g1932(.dina(\in1[122] ), .dinb(n2573), .dout(n2574));
  jor  g1933(.dina(n2574), .dinb(n2572), .dout(n2575));
  jnot g1934(.din(\in0[121] ), .dout(n2576));
  jand g1935(.dina(\in1[121] ), .dinb(n2576), .dout(n2577));
  jnot g1936(.din(\in0[120] ), .dout(n2578));
  jand g1937(.dina(\in1[120] ), .dinb(n2578), .dout(n2579));
  jor  g1938(.dina(n2579), .dinb(n2577), .dout(n2580));
  jor  g1939(.dina(n2580), .dinb(n2575), .dout(n2581));
  jnot g1940(.din(n2581), .dout(n2582));
  jand g1941(.dina(n2582), .dinb(n2570), .dout(n2583));
  jnot g1942(.din(\in1[123] ), .dout(n2584));
  jand g1943(.dina(n2584), .dinb(\in0[123] ), .dout(n2585));
  jnot g1944(.din(n2575), .dout(n2586));
  jnot g1945(.din(n2577), .dout(n2587));
  jnot g1946(.din(\in1[120] ), .dout(n2588));
  jand g1947(.dina(n2588), .dinb(\in0[120] ), .dout(n2589));
  jand g1948(.dina(n2589), .dinb(n2587), .dout(n2590));
  jnot g1949(.din(\in1[121] ), .dout(n2591));
  jand g1950(.dina(n2591), .dinb(\in0[121] ), .dout(n2592));
  jnot g1951(.din(\in1[122] ), .dout(n2593));
  jand g1952(.dina(n2593), .dinb(\in0[122] ), .dout(n2594));
  jor  g1953(.dina(n2594), .dinb(n2592), .dout(n2595));
  jor  g1954(.dina(n2595), .dinb(n2590), .dout(n2596));
  jand g1955(.dina(n2596), .dinb(n2586), .dout(n2597));
  jor  g1956(.dina(n2597), .dinb(n2585), .dout(n2598));
  jor  g1957(.dina(n2598), .dinb(n2583), .dout(n2599));
  jnot g1958(.din(\in0[126] ), .dout(n2600));
  jand g1959(.dina(\in1[126] ), .dinb(n2600), .dout(n2601));
  jnot g1960(.din(\in0[125] ), .dout(n2602));
  jand g1961(.dina(\in1[125] ), .dinb(n2602), .dout(n2603));
  jor  g1962(.dina(n2603), .dinb(n2601), .dout(n2604));
  jnot g1963(.din(\in1[127] ), .dout(n2605));
  jand g1964(.dina(n2605), .dinb(\in0[127] ), .dout(n2606));
  jnot g1965(.din(\in0[124] ), .dout(n2607));
  jand g1966(.dina(\in1[124] ), .dinb(n2607), .dout(n2608));
  jor  g1967(.dina(n2608), .dinb(n2606), .dout(n2609));
  jor  g1968(.dina(n2609), .dinb(n2604), .dout(n2610));
  jnot g1969(.din(n2610), .dout(n2611));
  jand g1970(.dina(n2611), .dinb(n2599), .dout(n2612));
  jnot g1971(.din(n2606), .dout(n2613));
  jnot g1972(.din(n2604), .dout(n2614));
  jnot g1973(.din(\in1[124] ), .dout(n2615));
  jand g1974(.dina(n2615), .dinb(\in0[124] ), .dout(n2616));
  jnot g1975(.din(\in1[125] ), .dout(n2617));
  jand g1976(.dina(n2617), .dinb(\in0[125] ), .dout(n2618));
  jor  g1977(.dina(n2618), .dinb(n2616), .dout(n2619));
  jand g1978(.dina(n2619), .dinb(n2614), .dout(n2620));
  jnot g1979(.din(\in1[126] ), .dout(n2621));
  jand g1980(.dina(n2621), .dinb(\in0[126] ), .dout(n2622));
  jor  g1981(.dina(n2622), .dinb(n2620), .dout(n2623));
  jand g1982(.dina(n2623), .dinb(n2613), .dout(n2624));
  jnot g1983(.din(\in0[127] ), .dout(n2625));
  jand g1984(.dina(\in1[127] ), .dinb(n2625), .dout(n2626));
  jor  g1985(.dina(n2626), .dinb(n2624), .dout(n2627));
  jor  g1986(.dina(n2627), .dinb(n2612), .dout(n2628));
  jand g1987(.dina(n2628), .dinb(\in0[30] ), .dout(n2629));
  jnot g1988(.din(n1718), .dout(n2630));
  jnot g1989(.din(n1723), .dout(n2631));
  jnot g1990(.din(n1728), .dout(n2632));
  jnot g1991(.din(n1733), .dout(n2633));
  jnot g1992(.din(n1738), .dout(n2634));
  jnot g1993(.din(n1743), .dout(n2635));
  jnot g1994(.din(n1748), .dout(n2636));
  jnot g1995(.din(n1753), .dout(n2637));
  jnot g1996(.din(n1758), .dout(n2638));
  jnot g1997(.din(n1763), .dout(n2639));
  jnot g1998(.din(n1768), .dout(n2640));
  jnot g1999(.din(n1773), .dout(n2641));
  jnot g2000(.din(n1778), .dout(n2642));
  jnot g2001(.din(n1783), .dout(n2643));
  jnot g2002(.din(n1788), .dout(n2644));
  jnot g2003(.din(n1793), .dout(n2645));
  jnot g2004(.din(n1798), .dout(n2646));
  jnot g2005(.din(n1803), .dout(n2647));
  jnot g2006(.din(n1808), .dout(n2648));
  jnot g2007(.din(n1813), .dout(n2649));
  jnot g2008(.din(n1818), .dout(n2650));
  jnot g2009(.din(n1823), .dout(n2651));
  jnot g2010(.din(n1828), .dout(n2652));
  jnot g2011(.din(n1833), .dout(n2653));
  jnot g2012(.din(n1838), .dout(n2654));
  jnot g2013(.din(n1843), .dout(n2655));
  jnot g2014(.din(n1848), .dout(n2656));
  jnot g2015(.din(n1853), .dout(n2657));
  jnot g2016(.din(\in0[1] ), .dout(n2658));
  jor  g2017(.dina(\in1[1] ), .dinb(n2658), .dout(n2659));
  jand g2018(.dina(\in1[1] ), .dinb(n2658), .dout(n2660));
  jnot g2019(.din(\in0[0] ), .dout(n2661));
  jor  g2020(.dina(\in1[0] ), .dinb(n2661), .dout(n2662));
  jor  g2021(.dina(n2662), .dinb(n2660), .dout(n2663));
  jand g2022(.dina(n2663), .dinb(n2659), .dout(n2664));
  jor  g2023(.dina(n2664), .dinb(n1855), .dout(n2665));
  jand g2024(.dina(n2665), .dinb(n2657), .dout(n2666));
  jor  g2025(.dina(n2666), .dinb(n1850), .dout(n2667));
  jand g2026(.dina(n2667), .dinb(n2656), .dout(n2668));
  jor  g2027(.dina(n2668), .dinb(n1845), .dout(n2669));
  jand g2028(.dina(n2669), .dinb(n2655), .dout(n2670));
  jor  g2029(.dina(n2670), .dinb(n1840), .dout(n2671));
  jand g2030(.dina(n2671), .dinb(n2654), .dout(n2672));
  jor  g2031(.dina(n2672), .dinb(n1835), .dout(n2673));
  jand g2032(.dina(n2673), .dinb(n2653), .dout(n2674));
  jor  g2033(.dina(n2674), .dinb(n1830), .dout(n2675));
  jand g2034(.dina(n2675), .dinb(n2652), .dout(n2676));
  jor  g2035(.dina(n2676), .dinb(n1825), .dout(n2677));
  jand g2036(.dina(n2677), .dinb(n2651), .dout(n2678));
  jor  g2037(.dina(n2678), .dinb(n1820), .dout(n2679));
  jand g2038(.dina(n2679), .dinb(n2650), .dout(n2680));
  jor  g2039(.dina(n2680), .dinb(n1815), .dout(n2681));
  jand g2040(.dina(n2681), .dinb(n2649), .dout(n2682));
  jor  g2041(.dina(n2682), .dinb(n1810), .dout(n2683));
  jand g2042(.dina(n2683), .dinb(n2648), .dout(n2684));
  jor  g2043(.dina(n2684), .dinb(n1805), .dout(n2685));
  jand g2044(.dina(n2685), .dinb(n2647), .dout(n2686));
  jor  g2045(.dina(n2686), .dinb(n1800), .dout(n2687));
  jand g2046(.dina(n2687), .dinb(n2646), .dout(n2688));
  jor  g2047(.dina(n2688), .dinb(n1795), .dout(n2689));
  jand g2048(.dina(n2689), .dinb(n2645), .dout(n2690));
  jor  g2049(.dina(n2690), .dinb(n1790), .dout(n2691));
  jand g2050(.dina(n2691), .dinb(n2644), .dout(n2692));
  jor  g2051(.dina(n2692), .dinb(n1785), .dout(n2693));
  jand g2052(.dina(n2693), .dinb(n2643), .dout(n2694));
  jor  g2053(.dina(n2694), .dinb(n1780), .dout(n2695));
  jand g2054(.dina(n2695), .dinb(n2642), .dout(n2696));
  jor  g2055(.dina(n2696), .dinb(n1775), .dout(n2697));
  jand g2056(.dina(n2697), .dinb(n2641), .dout(n2698));
  jor  g2057(.dina(n2698), .dinb(n1770), .dout(n2699));
  jand g2058(.dina(n2699), .dinb(n2640), .dout(n2700));
  jor  g2059(.dina(n2700), .dinb(n1765), .dout(n2701));
  jand g2060(.dina(n2701), .dinb(n2639), .dout(n2702));
  jor  g2061(.dina(n2702), .dinb(n1760), .dout(n2703));
  jand g2062(.dina(n2703), .dinb(n2638), .dout(n2704));
  jor  g2063(.dina(n2704), .dinb(n1755), .dout(n2705));
  jand g2064(.dina(n2705), .dinb(n2637), .dout(n2706));
  jor  g2065(.dina(n2706), .dinb(n1750), .dout(n2707));
  jand g2066(.dina(n2707), .dinb(n2636), .dout(n2708));
  jor  g2067(.dina(n2708), .dinb(n1745), .dout(n2709));
  jand g2068(.dina(n2709), .dinb(n2635), .dout(n2710));
  jor  g2069(.dina(n2710), .dinb(n1740), .dout(n2711));
  jand g2070(.dina(n2711), .dinb(n2634), .dout(n2712));
  jor  g2071(.dina(n2712), .dinb(n1735), .dout(n2713));
  jand g2072(.dina(n2713), .dinb(n2633), .dout(n2714));
  jor  g2073(.dina(n2714), .dinb(n1730), .dout(n2715));
  jand g2074(.dina(n2715), .dinb(n2632), .dout(n2716));
  jor  g2075(.dina(n2716), .dinb(n1725), .dout(n2717));
  jand g2076(.dina(n2717), .dinb(n2631), .dout(n2718));
  jor  g2077(.dina(n2718), .dinb(n1720), .dout(n2719));
  jand g2078(.dina(n2719), .dinb(n2630), .dout(n2720));
  jor  g2079(.dina(n2720), .dinb(n1715), .dout(n2721));
  jnot g2080(.din(n1925), .dout(n2722));
  jand g2081(.dina(n2722), .dinb(n2721), .dout(n2723));
  jor  g2082(.dina(n1952), .dinb(n2723), .dout(n2724));
  jnot g2083(.din(n1987), .dout(n2725));
  jand g2084(.dina(n2725), .dinb(n2724), .dout(n2726));
  jor  g2085(.dina(n2011), .dinb(n2726), .dout(n2727));
  jnot g2086(.din(n2046), .dout(n2728));
  jand g2087(.dina(n2728), .dinb(n2727), .dout(n2729));
  jor  g2088(.dina(n2073), .dinb(n2729), .dout(n2730));
  jnot g2089(.din(n2104), .dout(n2731));
  jand g2090(.dina(n2731), .dinb(n2730), .dout(n2732));
  jor  g2091(.dina(n2128), .dinb(n2732), .dout(n2733));
  jnot g2092(.din(n2163), .dout(n2734));
  jand g2093(.dina(n2734), .dinb(n2733), .dout(n2735));
  jor  g2094(.dina(n2175), .dinb(n2735), .dout(n2736));
  jnot g2095(.din(n2192), .dout(n2737));
  jand g2096(.dina(n2737), .dinb(n2736), .dout(n2738));
  jor  g2097(.dina(n2204), .dinb(n2738), .dout(n2739));
  jnot g2098(.din(n2221), .dout(n2740));
  jand g2099(.dina(n2740), .dinb(n2739), .dout(n2741));
  jor  g2100(.dina(n2233), .dinb(n2741), .dout(n2742));
  jnot g2101(.din(n2250), .dout(n2743));
  jand g2102(.dina(n2743), .dinb(n2742), .dout(n2744));
  jor  g2103(.dina(n2262), .dinb(n2744), .dout(n2745));
  jnot g2104(.din(n2279), .dout(n2746));
  jand g2105(.dina(n2746), .dinb(n2745), .dout(n2747));
  jor  g2106(.dina(n2291), .dinb(n2747), .dout(n2748));
  jnot g2107(.din(n2308), .dout(n2749));
  jand g2108(.dina(n2749), .dinb(n2748), .dout(n2750));
  jor  g2109(.dina(n2320), .dinb(n2750), .dout(n2751));
  jnot g2110(.din(n2337), .dout(n2752));
  jand g2111(.dina(n2752), .dinb(n2751), .dout(n2753));
  jor  g2112(.dina(n2349), .dinb(n2753), .dout(n2754));
  jnot g2113(.din(n2366), .dout(n2755));
  jand g2114(.dina(n2755), .dinb(n2754), .dout(n2756));
  jor  g2115(.dina(n2378), .dinb(n2756), .dout(n2757));
  jnot g2116(.din(n2395), .dout(n2758));
  jand g2117(.dina(n2758), .dinb(n2757), .dout(n2759));
  jor  g2118(.dina(n2407), .dinb(n2759), .dout(n2760));
  jnot g2119(.din(n2424), .dout(n2761));
  jand g2120(.dina(n2761), .dinb(n2760), .dout(n2762));
  jor  g2121(.dina(n2436), .dinb(n2762), .dout(n2763));
  jnot g2122(.din(n2453), .dout(n2764));
  jand g2123(.dina(n2764), .dinb(n2763), .dout(n2765));
  jor  g2124(.dina(n2465), .dinb(n2765), .dout(n2766));
  jnot g2125(.din(n2482), .dout(n2767));
  jand g2126(.dina(n2767), .dinb(n2766), .dout(n2768));
  jor  g2127(.dina(n2494), .dinb(n2768), .dout(n2769));
  jnot g2128(.din(n2511), .dout(n2770));
  jand g2129(.dina(n2770), .dinb(n2769), .dout(n2771));
  jor  g2130(.dina(n2523), .dinb(n2771), .dout(n2772));
  jnot g2131(.din(n2540), .dout(n2773));
  jand g2132(.dina(n2773), .dinb(n2772), .dout(n2774));
  jor  g2133(.dina(n2552), .dinb(n2774), .dout(n2775));
  jnot g2134(.din(n2569), .dout(n2776));
  jand g2135(.dina(n2776), .dinb(n2775), .dout(n2777));
  jor  g2136(.dina(n2581), .dinb(n2777), .dout(n2778));
  jnot g2137(.din(n2598), .dout(n2779));
  jand g2138(.dina(n2779), .dinb(n2778), .dout(n2780));
  jor  g2139(.dina(n2610), .dinb(n2780), .dout(n2781));
  jnot g2140(.din(n2627), .dout(n2782));
  jand g2141(.dina(n2782), .dinb(n2781), .dout(n2783));
  jand g2142(.dina(n2783), .dinb(\in1[30] ), .dout(n2784));
  jor  g2143(.dina(n2784), .dinb(n2629), .dout(n2785));
  jnot g2144(.din(n2785), .dout(n2786));
  jand g2145(.dina(n1556), .dinb(\in2[30] ), .dout(n2787));
  jand g2146(.dina(n1711), .dinb(\in3[30] ), .dout(n2788));
  jor  g2147(.dina(n2788), .dinb(n2787), .dout(n2789));
  jand g2148(.dina(n2789), .dinb(n2786), .dout(n2790));
  jand g2149(.dina(n2628), .dinb(\in0[29] ), .dout(n2791));
  jand g2150(.dina(n2783), .dinb(\in1[29] ), .dout(n2792));
  jor  g2151(.dina(n2792), .dinb(n2791), .dout(n2793));
  jand g2152(.dina(n1556), .dinb(\in2[29] ), .dout(n2794));
  jand g2153(.dina(n1711), .dinb(\in3[29] ), .dout(n2795));
  jor  g2154(.dina(n2795), .dinb(n2794), .dout(n2796));
  jnot g2155(.din(n2796), .dout(n2797));
  jand g2156(.dina(n2797), .dinb(n2793), .dout(n2798));
  jnot g2157(.din(n2798), .dout(n2799));
  jor  g2158(.dina(n2797), .dinb(n2793), .dout(n2800));
  jnot g2159(.din(n2800), .dout(n2801));
  jand g2160(.dina(n2628), .dinb(\in0[28] ), .dout(n2802));
  jand g2161(.dina(n2783), .dinb(\in1[28] ), .dout(n2803));
  jor  g2162(.dina(n2803), .dinb(n2802), .dout(n2804));
  jand g2163(.dina(n1556), .dinb(\in2[28] ), .dout(n2805));
  jand g2164(.dina(n1711), .dinb(\in3[28] ), .dout(n2806));
  jor  g2165(.dina(n2806), .dinb(n2805), .dout(n2807));
  jnot g2166(.din(n2807), .dout(n2808));
  jand g2167(.dina(n2808), .dinb(n2804), .dout(n2809));
  jnot g2168(.din(n2809), .dout(n2810));
  jor  g2169(.dina(n2808), .dinb(n2804), .dout(n2811));
  jnot g2170(.din(n2811), .dout(n2812));
  jand g2171(.dina(n2628), .dinb(\in0[27] ), .dout(n2813));
  jand g2172(.dina(n2783), .dinb(\in1[27] ), .dout(n2814));
  jor  g2173(.dina(n2814), .dinb(n2813), .dout(n2815));
  jand g2174(.dina(n1556), .dinb(\in2[27] ), .dout(n2816));
  jand g2175(.dina(n1711), .dinb(\in3[27] ), .dout(n2817));
  jor  g2176(.dina(n2817), .dinb(n2816), .dout(n2818));
  jnot g2177(.din(n2818), .dout(n2819));
  jand g2178(.dina(n2819), .dinb(n2815), .dout(n2820));
  jnot g2179(.din(n2820), .dout(n2821));
  jor  g2180(.dina(n2819), .dinb(n2815), .dout(n2822));
  jnot g2181(.din(n2822), .dout(n2823));
  jand g2182(.dina(n2628), .dinb(\in0[26] ), .dout(n2824));
  jand g2183(.dina(n2783), .dinb(\in1[26] ), .dout(n2825));
  jor  g2184(.dina(n2825), .dinb(n2824), .dout(n2826));
  jand g2185(.dina(n1556), .dinb(\in2[26] ), .dout(n2827));
  jand g2186(.dina(n1711), .dinb(\in3[26] ), .dout(n2828));
  jor  g2187(.dina(n2828), .dinb(n2827), .dout(n2829));
  jnot g2188(.din(n2829), .dout(n2830));
  jand g2189(.dina(n2830), .dinb(n2826), .dout(n2831));
  jnot g2190(.din(n2831), .dout(n2832));
  jor  g2191(.dina(n2830), .dinb(n2826), .dout(n2833));
  jnot g2192(.din(n2833), .dout(n2834));
  jand g2193(.dina(n2628), .dinb(\in0[25] ), .dout(n2835));
  jand g2194(.dina(n2783), .dinb(\in1[25] ), .dout(n2836));
  jor  g2195(.dina(n2836), .dinb(n2835), .dout(n2837));
  jand g2196(.dina(n1556), .dinb(\in2[25] ), .dout(n2838));
  jand g2197(.dina(n1711), .dinb(\in3[25] ), .dout(n2839));
  jor  g2198(.dina(n2839), .dinb(n2838), .dout(n2840));
  jnot g2199(.din(n2840), .dout(n2841));
  jand g2200(.dina(n2841), .dinb(n2837), .dout(n2842));
  jnot g2201(.din(n2842), .dout(n2843));
  jor  g2202(.dina(n2841), .dinb(n2837), .dout(n2844));
  jnot g2203(.din(n2844), .dout(n2845));
  jand g2204(.dina(n2628), .dinb(\in0[24] ), .dout(n2846));
  jand g2205(.dina(n2783), .dinb(\in1[24] ), .dout(n2847));
  jor  g2206(.dina(n2847), .dinb(n2846), .dout(n2848));
  jand g2207(.dina(n1556), .dinb(\in2[24] ), .dout(n2849));
  jand g2208(.dina(n1711), .dinb(\in3[24] ), .dout(n2850));
  jor  g2209(.dina(n2850), .dinb(n2849), .dout(n2851));
  jnot g2210(.din(n2851), .dout(n2852));
  jand g2211(.dina(n2852), .dinb(n2848), .dout(n2853));
  jnot g2212(.din(n2853), .dout(n2854));
  jand g2213(.dina(n2628), .dinb(\in0[22] ), .dout(n2855));
  jand g2214(.dina(n2783), .dinb(\in1[22] ), .dout(n2856));
  jor  g2215(.dina(n2856), .dinb(n2855), .dout(n2857));
  jnot g2216(.din(n2857), .dout(n2858));
  jand g2217(.dina(n1556), .dinb(\in2[22] ), .dout(n2859));
  jand g2218(.dina(n1711), .dinb(\in3[22] ), .dout(n2860));
  jor  g2219(.dina(n2860), .dinb(n2859), .dout(n2861));
  jand g2220(.dina(n2861), .dinb(n2858), .dout(n2862));
  jand g2221(.dina(n2628), .dinb(\in0[21] ), .dout(n2863));
  jand g2222(.dina(n2783), .dinb(\in1[21] ), .dout(n2864));
  jor  g2223(.dina(n2864), .dinb(n2863), .dout(n2865));
  jand g2224(.dina(n1556), .dinb(\in2[21] ), .dout(n2866));
  jand g2225(.dina(n1711), .dinb(\in3[21] ), .dout(n2867));
  jor  g2226(.dina(n2867), .dinb(n2866), .dout(n2868));
  jnot g2227(.din(n2868), .dout(n2869));
  jand g2228(.dina(n2869), .dinb(n2865), .dout(n2870));
  jnot g2229(.din(n2870), .dout(n2871));
  jor  g2230(.dina(n2869), .dinb(n2865), .dout(n2872));
  jnot g2231(.din(n2872), .dout(n2873));
  jand g2232(.dina(n2628), .dinb(\in0[20] ), .dout(n2874));
  jand g2233(.dina(n2783), .dinb(\in1[20] ), .dout(n2875));
  jor  g2234(.dina(n2875), .dinb(n2874), .dout(n2876));
  jand g2235(.dina(n1556), .dinb(\in2[20] ), .dout(n2877));
  jand g2236(.dina(n1711), .dinb(\in3[20] ), .dout(n2878));
  jor  g2237(.dina(n2878), .dinb(n2877), .dout(n2879));
  jnot g2238(.din(n2879), .dout(n2880));
  jand g2239(.dina(n2880), .dinb(n2876), .dout(n2881));
  jnot g2240(.din(n2881), .dout(n2882));
  jor  g2241(.dina(n2880), .dinb(n2876), .dout(n2883));
  jnot g2242(.din(n2883), .dout(n2884));
  jand g2243(.dina(n2628), .dinb(\in0[19] ), .dout(n2885));
  jand g2244(.dina(n2783), .dinb(\in1[19] ), .dout(n2886));
  jor  g2245(.dina(n2886), .dinb(n2885), .dout(n2887));
  jand g2246(.dina(n1556), .dinb(\in2[19] ), .dout(n2888));
  jand g2247(.dina(n1711), .dinb(\in3[19] ), .dout(n2889));
  jor  g2248(.dina(n2889), .dinb(n2888), .dout(n2890));
  jnot g2249(.din(n2890), .dout(n2891));
  jand g2250(.dina(n2891), .dinb(n2887), .dout(n2892));
  jnot g2251(.din(n2892), .dout(n2893));
  jand g2252(.dina(n1556), .dinb(\in2[17] ), .dout(n2894));
  jand g2253(.dina(n1711), .dinb(\in3[17] ), .dout(n2895));
  jor  g2254(.dina(n2895), .dinb(n2894), .dout(n2896));
  jand g2255(.dina(n2628), .dinb(\in0[17] ), .dout(n2897));
  jand g2256(.dina(n2783), .dinb(\in1[17] ), .dout(n2898));
  jor  g2257(.dina(n2898), .dinb(n2897), .dout(n2899));
  jnot g2258(.din(n2899), .dout(n2900));
  jand g2259(.dina(n2628), .dinb(\in0[16] ), .dout(n2901));
  jand g2260(.dina(n2783), .dinb(\in1[16] ), .dout(n2902));
  jor  g2261(.dina(n2902), .dinb(n2901), .dout(n2903));
  jnot g2262(.din(n2903), .dout(n2904));
  jand g2263(.dina(n1556), .dinb(\in2[16] ), .dout(n2905));
  jand g2264(.dina(n1711), .dinb(\in3[16] ), .dout(n2906));
  jor  g2265(.dina(n2906), .dinb(n2905), .dout(n2907));
  jand g2266(.dina(n2907), .dinb(n2904), .dout(n2908));
  jor  g2267(.dina(n2907), .dinb(n2904), .dout(n2909));
  jand g2268(.dina(n2628), .dinb(\in0[15] ), .dout(n2910));
  jand g2269(.dina(n2783), .dinb(\in1[15] ), .dout(n2911));
  jor  g2270(.dina(n2911), .dinb(n2910), .dout(n2912));
  jnot g2271(.din(n2912), .dout(n2913));
  jand g2272(.dina(n1556), .dinb(\in2[15] ), .dout(n2914));
  jand g2273(.dina(n1711), .dinb(\in3[15] ), .dout(n2915));
  jor  g2274(.dina(n2915), .dinb(n2914), .dout(n2916));
  jand g2275(.dina(n2916), .dinb(n2913), .dout(n2917));
  jand g2276(.dina(n2628), .dinb(\in0[14] ), .dout(n2918));
  jand g2277(.dina(n2783), .dinb(\in1[14] ), .dout(n2919));
  jor  g2278(.dina(n2919), .dinb(n2918), .dout(n2920));
  jnot g2279(.din(n2920), .dout(n2921));
  jand g2280(.dina(n1556), .dinb(\in2[14] ), .dout(n2922));
  jand g2281(.dina(n1711), .dinb(\in3[14] ), .dout(n2923));
  jor  g2282(.dina(n2923), .dinb(n2922), .dout(n2924));
  jand g2283(.dina(n2924), .dinb(n2921), .dout(n2925));
  jand g2284(.dina(n2628), .dinb(\in0[13] ), .dout(n2926));
  jand g2285(.dina(n2783), .dinb(\in1[13] ), .dout(n2927));
  jor  g2286(.dina(n2927), .dinb(n2926), .dout(n2928));
  jand g2287(.dina(n1556), .dinb(\in2[13] ), .dout(n2929));
  jand g2288(.dina(n1711), .dinb(\in3[13] ), .dout(n2930));
  jor  g2289(.dina(n2930), .dinb(n2929), .dout(n2931));
  jnot g2290(.din(n2931), .dout(n2932));
  jand g2291(.dina(n2932), .dinb(n2928), .dout(n2933));
  jnot g2292(.din(n2933), .dout(n2934));
  jor  g2293(.dina(n2932), .dinb(n2928), .dout(n2935));
  jnot g2294(.din(n2935), .dout(n2936));
  jand g2295(.dina(n2628), .dinb(\in0[12] ), .dout(n2937));
  jand g2296(.dina(n2783), .dinb(\in1[12] ), .dout(n2938));
  jor  g2297(.dina(n2938), .dinb(n2937), .dout(n2939));
  jand g2298(.dina(n1556), .dinb(\in2[12] ), .dout(n2940));
  jand g2299(.dina(n1711), .dinb(\in3[12] ), .dout(n2941));
  jor  g2300(.dina(n2941), .dinb(n2940), .dout(n2942));
  jnot g2301(.din(n2942), .dout(n2943));
  jand g2302(.dina(n2943), .dinb(n2939), .dout(n2944));
  jnot g2303(.din(n2944), .dout(n2945));
  jor  g2304(.dina(n2943), .dinb(n2939), .dout(n2946));
  jnot g2305(.din(n2946), .dout(n2947));
  jand g2306(.dina(n2628), .dinb(\in0[11] ), .dout(n2948));
  jand g2307(.dina(n2783), .dinb(\in1[11] ), .dout(n2949));
  jor  g2308(.dina(n2949), .dinb(n2948), .dout(n2950));
  jand g2309(.dina(n1556), .dinb(\in2[11] ), .dout(n2951));
  jand g2310(.dina(n1711), .dinb(\in3[11] ), .dout(n2952));
  jor  g2311(.dina(n2952), .dinb(n2951), .dout(n2953));
  jnot g2312(.din(n2953), .dout(n2954));
  jand g2313(.dina(n2954), .dinb(n2950), .dout(n2955));
  jnot g2314(.din(n2955), .dout(n2956));
  jor  g2315(.dina(n2954), .dinb(n2950), .dout(n2957));
  jnot g2316(.din(n2957), .dout(n2958));
  jand g2317(.dina(n2628), .dinb(\in0[10] ), .dout(n2959));
  jand g2318(.dina(n2783), .dinb(\in1[10] ), .dout(n2960));
  jor  g2319(.dina(n2960), .dinb(n2959), .dout(n2961));
  jand g2320(.dina(n1556), .dinb(\in2[10] ), .dout(n2962));
  jand g2321(.dina(n1711), .dinb(\in3[10] ), .dout(n2963));
  jor  g2322(.dina(n2963), .dinb(n2962), .dout(n2964));
  jnot g2323(.din(n2964), .dout(n2965));
  jand g2324(.dina(n2965), .dinb(n2961), .dout(n2966));
  jnot g2325(.din(n2966), .dout(n2967));
  jor  g2326(.dina(n2965), .dinb(n2961), .dout(n2968));
  jnot g2327(.din(n2968), .dout(n2969));
  jand g2328(.dina(n2628), .dinb(\in0[9] ), .dout(n2970));
  jand g2329(.dina(n2783), .dinb(\in1[9] ), .dout(n2971));
  jor  g2330(.dina(n2971), .dinb(n2970), .dout(n2972));
  jand g2331(.dina(n1556), .dinb(\in2[9] ), .dout(n2973));
  jand g2332(.dina(n1711), .dinb(\in3[9] ), .dout(n2974));
  jor  g2333(.dina(n2974), .dinb(n2973), .dout(n2975));
  jnot g2334(.din(n2975), .dout(n2976));
  jand g2335(.dina(n2976), .dinb(n2972), .dout(n2977));
  jnot g2336(.din(n2977), .dout(n2978));
  jor  g2337(.dina(n2976), .dinb(n2972), .dout(n2979));
  jnot g2338(.din(n2979), .dout(n2980));
  jand g2339(.dina(n1556), .dinb(\in2[8] ), .dout(n2981));
  jand g2340(.dina(n1711), .dinb(\in3[8] ), .dout(n2982));
  jor  g2341(.dina(n2982), .dinb(n2981), .dout(n2983));
  jand g2342(.dina(n2628), .dinb(\in0[7] ), .dout(n2984));
  jand g2343(.dina(n2783), .dinb(\in1[7] ), .dout(n2985));
  jor  g2344(.dina(n2985), .dinb(n2984), .dout(n2986));
  jand g2345(.dina(n1556), .dinb(\in2[7] ), .dout(n2987));
  jand g2346(.dina(n1711), .dinb(\in3[7] ), .dout(n2988));
  jor  g2347(.dina(n2988), .dinb(n2987), .dout(n2989));
  jnot g2348(.din(n2989), .dout(n2990));
  jand g2349(.dina(n2990), .dinb(n2986), .dout(n2991));
  jnot g2350(.din(n2991), .dout(n2992));
  jor  g2351(.dina(n2990), .dinb(n2986), .dout(n2993));
  jnot g2352(.din(n2993), .dout(n2994));
  jand g2353(.dina(n2628), .dinb(\in0[5] ), .dout(n2995));
  jand g2354(.dina(n2783), .dinb(\in1[5] ), .dout(n2996));
  jor  g2355(.dina(n2996), .dinb(n2995), .dout(n2997));
  jnot g2356(.din(n2997), .dout(n2998));
  jand g2357(.dina(n2628), .dinb(\in0[4] ), .dout(n2999));
  jand g2358(.dina(n2783), .dinb(\in1[4] ), .dout(n3000));
  jor  g2359(.dina(n3000), .dinb(n2999), .dout(n3001));
  jnot g2360(.din(n3001), .dout(n3002));
  jand g2361(.dina(n2628), .dinb(\in0[3] ), .dout(n3003));
  jand g2362(.dina(n2783), .dinb(\in1[3] ), .dout(n3004));
  jor  g2363(.dina(n3004), .dinb(n3003), .dout(n3005));
  jnot g2364(.din(n3005), .dout(n3006));
  jand g2365(.dina(n1556), .dinb(\in2[3] ), .dout(n3007));
  jand g2366(.dina(n1711), .dinb(\in3[3] ), .dout(n3008));
  jor  g2367(.dina(n3008), .dinb(n3007), .dout(n3009));
  jand g2368(.dina(n3009), .dinb(n3006), .dout(n3010));
  jor  g2369(.dina(n3009), .dinb(n3006), .dout(n3011));
  jor  g2370(.dina(n2783), .dinb(n1854), .dout(n3012));
  jor  g2371(.dina(n2628), .dinb(n1852), .dout(n3013));
  jand g2372(.dina(n3013), .dinb(n3012), .dout(n3014));
  jand g2373(.dina(n1556), .dinb(\in2[2] ), .dout(n3015));
  jand g2374(.dina(n1711), .dinb(\in3[2] ), .dout(n3016));
  jor  g2375(.dina(n3016), .dinb(n3015), .dout(n3017));
  jand g2376(.dina(n3017), .dinb(n3014), .dout(n3018));
  jand g2377(.dina(n1556), .dinb(\in2[1] ), .dout(n3019));
  jand g2378(.dina(n1711), .dinb(\in3[1] ), .dout(n3020));
  jor  g2379(.dina(n3020), .dinb(n3019), .dout(n3021));
  jor  g2380(.dina(n2783), .dinb(n2661), .dout(n3022));
  jor  g2381(.dina(n2628), .dinb(n1860), .dout(n3023));
  jand g2382(.dina(n3023), .dinb(n3022), .dout(n3024));
  jor  g2383(.dina(n3024), .dinb(n1713), .dout(n3025));
  jor  g2384(.dina(n2783), .dinb(n2658), .dout(n3026));
  jor  g2385(.dina(n2628), .dinb(n1857), .dout(n3027));
  jand g2386(.dina(n3027), .dinb(n3026), .dout(n3028));
  jand g2387(.dina(n3028), .dinb(n3025), .dout(n3029));
  jor  g2388(.dina(n3029), .dinb(n3021), .dout(n3030));
  jor  g2389(.dina(n3017), .dinb(n3014), .dout(n3031));
  jor  g2390(.dina(n3028), .dinb(n3025), .dout(n3032));
  jand g2391(.dina(n3032), .dinb(n3031), .dout(n3033));
  jand g2392(.dina(n3033), .dinb(n3030), .dout(n3034));
  jor  g2393(.dina(n3034), .dinb(n3018), .dout(n3035));
  jand g2394(.dina(n3035), .dinb(n3011), .dout(n3036));
  jor  g2395(.dina(n3036), .dinb(n3010), .dout(n3037));
  jand g2396(.dina(n1556), .dinb(\in2[4] ), .dout(n3038));
  jand g2397(.dina(n1711), .dinb(\in3[4] ), .dout(n3039));
  jor  g2398(.dina(n3039), .dinb(n3038), .dout(n3040));
  jor  g2399(.dina(n3040), .dinb(n3037), .dout(n3041));
  jand g2400(.dina(n3041), .dinb(n3002), .dout(n3042));
  jand g2401(.dina(n3040), .dinb(n3037), .dout(n3043));
  jor  g2402(.dina(n3043), .dinb(n3042), .dout(n3044));
  jand g2403(.dina(n1556), .dinb(\in2[5] ), .dout(n3045));
  jand g2404(.dina(n1711), .dinb(\in3[5] ), .dout(n3046));
  jor  g2405(.dina(n3046), .dinb(n3045), .dout(n3047));
  jor  g2406(.dina(n3047), .dinb(n3044), .dout(n3048));
  jand g2407(.dina(n3048), .dinb(n2998), .dout(n3049));
  jand g2408(.dina(n3047), .dinb(n3044), .dout(n3050));
  jand g2409(.dina(n2628), .dinb(\in0[6] ), .dout(n3051));
  jand g2410(.dina(n2783), .dinb(\in1[6] ), .dout(n3052));
  jor  g2411(.dina(n3052), .dinb(n3051), .dout(n3053));
  jnot g2412(.din(n3053), .dout(n3054));
  jand g2413(.dina(n1556), .dinb(\in2[6] ), .dout(n3055));
  jand g2414(.dina(n1711), .dinb(\in3[6] ), .dout(n3056));
  jor  g2415(.dina(n3056), .dinb(n3055), .dout(n3057));
  jand g2416(.dina(n3057), .dinb(n3054), .dout(n3058));
  jor  g2417(.dina(n3058), .dinb(n3050), .dout(n3059));
  jor  g2418(.dina(n3059), .dinb(n3049), .dout(n3060));
  jor  g2419(.dina(n3057), .dinb(n3054), .dout(n3061));
  jand g2420(.dina(n3061), .dinb(n3060), .dout(n3062));
  jor  g2421(.dina(n3062), .dinb(n2994), .dout(n3063));
  jand g2422(.dina(n3063), .dinb(n2992), .dout(n3064));
  jand g2423(.dina(n2628), .dinb(\in0[8] ), .dout(n3065));
  jand g2424(.dina(n2783), .dinb(\in1[8] ), .dout(n3066));
  jor  g2425(.dina(n3066), .dinb(n3065), .dout(n3067));
  jnot g2426(.din(n3067), .dout(n3068));
  jand g2427(.dina(n3068), .dinb(n3064), .dout(n3069));
  jor  g2428(.dina(n3069), .dinb(n2983), .dout(n3070));
  jor  g2429(.dina(n3068), .dinb(n3064), .dout(n3071));
  jand g2430(.dina(n3071), .dinb(n3070), .dout(n3072));
  jor  g2431(.dina(n3072), .dinb(n2980), .dout(n3073));
  jand g2432(.dina(n3073), .dinb(n2978), .dout(n3074));
  jor  g2433(.dina(n3074), .dinb(n2969), .dout(n3075));
  jand g2434(.dina(n3075), .dinb(n2967), .dout(n3076));
  jor  g2435(.dina(n3076), .dinb(n2958), .dout(n3077));
  jand g2436(.dina(n3077), .dinb(n2956), .dout(n3078));
  jor  g2437(.dina(n3078), .dinb(n2947), .dout(n3079));
  jand g2438(.dina(n3079), .dinb(n2945), .dout(n3080));
  jor  g2439(.dina(n3080), .dinb(n2936), .dout(n3081));
  jand g2440(.dina(n3081), .dinb(n2934), .dout(n3082));
  jor  g2441(.dina(n3082), .dinb(n2925), .dout(n3083));
  jor  g2442(.dina(n2924), .dinb(n2921), .dout(n3084));
  jor  g2443(.dina(n2916), .dinb(n2913), .dout(n3085));
  jand g2444(.dina(n3085), .dinb(n3084), .dout(n3086));
  jand g2445(.dina(n3086), .dinb(n3083), .dout(n3087));
  jor  g2446(.dina(n3087), .dinb(n2917), .dout(n3088));
  jand g2447(.dina(n3088), .dinb(n2909), .dout(n3089));
  jor  g2448(.dina(n3089), .dinb(n2908), .dout(n3090));
  jand g2449(.dina(n3090), .dinb(n2900), .dout(n3091));
  jor  g2450(.dina(n3091), .dinb(n2896), .dout(n3092));
  jand g2451(.dina(n2628), .dinb(\in0[18] ), .dout(n3093));
  jand g2452(.dina(n2783), .dinb(\in1[18] ), .dout(n3094));
  jor  g2453(.dina(n3094), .dinb(n3093), .dout(n3095));
  jand g2454(.dina(n1556), .dinb(\in2[18] ), .dout(n3096));
  jand g2455(.dina(n1711), .dinb(\in3[18] ), .dout(n3097));
  jor  g2456(.dina(n3097), .dinb(n3096), .dout(n3098));
  jnot g2457(.din(n3098), .dout(n3099));
  jand g2458(.dina(n3099), .dinb(n3095), .dout(n3100));
  jnot g2459(.din(n3100), .dout(n3101));
  jor  g2460(.dina(n3090), .dinb(n2900), .dout(n3102));
  jand g2461(.dina(n3102), .dinb(n3101), .dout(n3103));
  jand g2462(.dina(n3103), .dinb(n3092), .dout(n3104));
  jor  g2463(.dina(n2891), .dinb(n2887), .dout(n3105));
  jor  g2464(.dina(n3099), .dinb(n3095), .dout(n3106));
  jand g2465(.dina(n3106), .dinb(n3105), .dout(n3107));
  jnot g2466(.din(n3107), .dout(n3108));
  jor  g2467(.dina(n3108), .dinb(n3104), .dout(n3109));
  jand g2468(.dina(n3109), .dinb(n2893), .dout(n3110));
  jor  g2469(.dina(n3110), .dinb(n2884), .dout(n3111));
  jand g2470(.dina(n3111), .dinb(n2882), .dout(n3112));
  jor  g2471(.dina(n3112), .dinb(n2873), .dout(n3113));
  jand g2472(.dina(n3113), .dinb(n2871), .dout(n3114));
  jor  g2473(.dina(n3114), .dinb(n2862), .dout(n3115));
  jor  g2474(.dina(n2861), .dinb(n2858), .dout(n3116));
  jand g2475(.dina(n2628), .dinb(\in0[23] ), .dout(n3117));
  jand g2476(.dina(n2783), .dinb(\in1[23] ), .dout(n3118));
  jor  g2477(.dina(n3118), .dinb(n3117), .dout(n3119));
  jand g2478(.dina(n1556), .dinb(\in2[23] ), .dout(n3120));
  jand g2479(.dina(n1711), .dinb(\in3[23] ), .dout(n3121));
  jor  g2480(.dina(n3121), .dinb(n3120), .dout(n3122));
  jnot g2481(.din(n3122), .dout(n3123));
  jand g2482(.dina(n3123), .dinb(n3119), .dout(n3124));
  jnot g2483(.din(n3124), .dout(n3125));
  jand g2484(.dina(n3125), .dinb(n3116), .dout(n3126));
  jand g2485(.dina(n3126), .dinb(n3115), .dout(n3127));
  jor  g2486(.dina(n3123), .dinb(n3119), .dout(n3128));
  jor  g2487(.dina(n2852), .dinb(n2848), .dout(n3129));
  jand g2488(.dina(n3129), .dinb(n3128), .dout(n3130));
  jnot g2489(.din(n3130), .dout(n3131));
  jor  g2490(.dina(n3131), .dinb(n3127), .dout(n3132));
  jand g2491(.dina(n3132), .dinb(n2854), .dout(n3133));
  jor  g2492(.dina(n3133), .dinb(n2845), .dout(n3134));
  jand g2493(.dina(n3134), .dinb(n2843), .dout(n3135));
  jor  g2494(.dina(n3135), .dinb(n2834), .dout(n3136));
  jand g2495(.dina(n3136), .dinb(n2832), .dout(n3137));
  jor  g2496(.dina(n3137), .dinb(n2823), .dout(n3138));
  jand g2497(.dina(n3138), .dinb(n2821), .dout(n3139));
  jor  g2498(.dina(n3139), .dinb(n2812), .dout(n3140));
  jand g2499(.dina(n3140), .dinb(n2810), .dout(n3141));
  jor  g2500(.dina(n3141), .dinb(n2801), .dout(n3142));
  jand g2501(.dina(n3142), .dinb(n2799), .dout(n3143));
  jor  g2502(.dina(n3143), .dinb(n2790), .dout(n3144));
  jor  g2503(.dina(n2789), .dinb(n2786), .dout(n3145));
  jand g2504(.dina(n2628), .dinb(\in0[31] ), .dout(n3146));
  jand g2505(.dina(n2783), .dinb(\in1[31] ), .dout(n3147));
  jor  g2506(.dina(n3147), .dinb(n3146), .dout(n3148));
  jand g2507(.dina(n1556), .dinb(\in2[31] ), .dout(n3149));
  jand g2508(.dina(n1711), .dinb(\in3[31] ), .dout(n3150));
  jor  g2509(.dina(n3150), .dinb(n3149), .dout(n3151));
  jnot g2510(.din(n3151), .dout(n3152));
  jand g2511(.dina(n3152), .dinb(n3148), .dout(n3153));
  jnot g2512(.din(n3153), .dout(n3154));
  jand g2513(.dina(n3154), .dinb(n3145), .dout(n3155));
  jand g2514(.dina(n3155), .dinb(n3144), .dout(n3156));
  jand g2515(.dina(n2628), .dinb(\in0[37] ), .dout(n3157));
  jand g2516(.dina(n2783), .dinb(\in1[37] ), .dout(n3158));
  jor  g2517(.dina(n3158), .dinb(n3157), .dout(n3159));
  jnot g2518(.din(n3159), .dout(n3160));
  jand g2519(.dina(n1556), .dinb(\in2[37] ), .dout(n3161));
  jand g2520(.dina(n1711), .dinb(\in3[37] ), .dout(n3162));
  jor  g2521(.dina(n3162), .dinb(n3161), .dout(n3163));
  jand g2522(.dina(n3163), .dinb(n3160), .dout(n3164));
  jand g2523(.dina(n2628), .dinb(\in0[39] ), .dout(n3165));
  jand g2524(.dina(n2783), .dinb(\in1[39] ), .dout(n3166));
  jor  g2525(.dina(n3166), .dinb(n3165), .dout(n3167));
  jnot g2526(.din(n3167), .dout(n3168));
  jand g2527(.dina(n1556), .dinb(\in2[39] ), .dout(n3169));
  jand g2528(.dina(n1711), .dinb(\in3[39] ), .dout(n3170));
  jor  g2529(.dina(n3170), .dinb(n3169), .dout(n3171));
  jand g2530(.dina(n3171), .dinb(n3168), .dout(n3172));
  jand g2531(.dina(n1556), .dinb(\in2[38] ), .dout(n3173));
  jand g2532(.dina(n1711), .dinb(\in3[38] ), .dout(n3174));
  jor  g2533(.dina(n3174), .dinb(n3173), .dout(n3175));
  jand g2534(.dina(n2628), .dinb(\in0[38] ), .dout(n3176));
  jand g2535(.dina(n2783), .dinb(\in1[38] ), .dout(n3177));
  jor  g2536(.dina(n3177), .dinb(n3176), .dout(n3178));
  jnot g2537(.din(n3178), .dout(n3179));
  jand g2538(.dina(n3179), .dinb(n3175), .dout(n3180));
  jor  g2539(.dina(n3180), .dinb(n3172), .dout(n3181));
  jor  g2540(.dina(n3181), .dinb(n3164), .dout(n3182));
  jnot g2541(.din(n3182), .dout(n3183));
  jand g2542(.dina(n2628), .dinb(\in0[35] ), .dout(n3184));
  jand g2543(.dina(n2783), .dinb(\in1[35] ), .dout(n3185));
  jor  g2544(.dina(n3185), .dinb(n3184), .dout(n3186));
  jnot g2545(.din(n3186), .dout(n3187));
  jand g2546(.dina(n1556), .dinb(\in2[35] ), .dout(n3188));
  jand g2547(.dina(n1711), .dinb(\in3[35] ), .dout(n3189));
  jor  g2548(.dina(n3189), .dinb(n3188), .dout(n3190));
  jand g2549(.dina(n3190), .dinb(n3187), .dout(n3191));
  jand g2550(.dina(n2628), .dinb(\in0[33] ), .dout(n3192));
  jand g2551(.dina(n2783), .dinb(\in1[33] ), .dout(n3193));
  jor  g2552(.dina(n3193), .dinb(n3192), .dout(n3194));
  jnot g2553(.din(n3194), .dout(n3195));
  jand g2554(.dina(n1556), .dinb(\in2[33] ), .dout(n3196));
  jand g2555(.dina(n1711), .dinb(\in3[33] ), .dout(n3197));
  jor  g2556(.dina(n3197), .dinb(n3196), .dout(n3198));
  jand g2557(.dina(n3198), .dinb(n3195), .dout(n3199));
  jand g2558(.dina(n1556), .dinb(\in2[34] ), .dout(n3200));
  jand g2559(.dina(n1711), .dinb(\in3[34] ), .dout(n3201));
  jor  g2560(.dina(n3201), .dinb(n3200), .dout(n3202));
  jand g2561(.dina(n2628), .dinb(\in0[34] ), .dout(n3203));
  jand g2562(.dina(n2783), .dinb(\in1[34] ), .dout(n3204));
  jor  g2563(.dina(n3204), .dinb(n3203), .dout(n3205));
  jnot g2564(.din(n3205), .dout(n3206));
  jand g2565(.dina(n3206), .dinb(n3202), .dout(n3207));
  jor  g2566(.dina(n3207), .dinb(n3199), .dout(n3208));
  jor  g2567(.dina(n3208), .dinb(n3191), .dout(n3209));
  jnot g2568(.din(n3209), .dout(n3210));
  jand g2569(.dina(n1556), .dinb(\in2[32] ), .dout(n3211));
  jand g2570(.dina(n1711), .dinb(\in3[32] ), .dout(n3212));
  jor  g2571(.dina(n3212), .dinb(n3211), .dout(n3213));
  jand g2572(.dina(n2628), .dinb(\in0[32] ), .dout(n3214));
  jand g2573(.dina(n2783), .dinb(\in1[32] ), .dout(n3215));
  jor  g2574(.dina(n3215), .dinb(n3214), .dout(n3216));
  jnot g2575(.din(n3216), .dout(n3217));
  jand g2576(.dina(n3217), .dinb(n3213), .dout(n3218));
  jnot g2577(.din(n3218), .dout(n3219));
  jand g2578(.dina(n2628), .dinb(\in0[36] ), .dout(n3220));
  jand g2579(.dina(n2783), .dinb(\in1[36] ), .dout(n3221));
  jor  g2580(.dina(n3221), .dinb(n3220), .dout(n3222));
  jnot g2581(.din(n3222), .dout(n3223));
  jand g2582(.dina(n1556), .dinb(\in2[36] ), .dout(n3224));
  jand g2583(.dina(n1711), .dinb(\in3[36] ), .dout(n3225));
  jor  g2584(.dina(n3225), .dinb(n3224), .dout(n3226));
  jand g2585(.dina(n3226), .dinb(n3223), .dout(n3227));
  jnot g2586(.din(n3227), .dout(n3228));
  jor  g2587(.dina(n3152), .dinb(n3148), .dout(n3229));
  jand g2588(.dina(n3229), .dinb(n3228), .dout(n3230));
  jand g2589(.dina(n3230), .dinb(n3219), .dout(n3231));
  jand g2590(.dina(n3231), .dinb(n3210), .dout(n3232));
  jand g2591(.dina(n3232), .dinb(n3183), .dout(n3233));
  jnot g2592(.din(n3233), .dout(n3234));
  jor  g2593(.dina(n3234), .dinb(n3156), .dout(n3235));
  jor  g2594(.dina(n3217), .dinb(n3213), .dout(n3236));
  jor  g2595(.dina(n3198), .dinb(n3195), .dout(n3237));
  jand g2596(.dina(n3237), .dinb(n3236), .dout(n3238));
  jor  g2597(.dina(n3238), .dinb(n3209), .dout(n3239));
  jor  g2598(.dina(n3206), .dinb(n3202), .dout(n3240));
  jor  g2599(.dina(n3240), .dinb(n3191), .dout(n3241));
  jor  g2600(.dina(n3190), .dinb(n3187), .dout(n3242));
  jand g2601(.dina(n3242), .dinb(n3241), .dout(n3243));
  jand g2602(.dina(n3243), .dinb(n3239), .dout(n3244));
  jor  g2603(.dina(n3244), .dinb(n3227), .dout(n3245));
  jor  g2604(.dina(n3226), .dinb(n3223), .dout(n3246));
  jor  g2605(.dina(n3163), .dinb(n3160), .dout(n3247));
  jand g2606(.dina(n3247), .dinb(n3246), .dout(n3248));
  jand g2607(.dina(n3248), .dinb(n3245), .dout(n3249));
  jor  g2608(.dina(n3249), .dinb(n3182), .dout(n3250));
  jor  g2609(.dina(n3179), .dinb(n3175), .dout(n3251));
  jor  g2610(.dina(n3251), .dinb(n3172), .dout(n3252));
  jor  g2611(.dina(n3171), .dinb(n3168), .dout(n3253));
  jand g2612(.dina(n3253), .dinb(n3252), .dout(n3254));
  jand g2613(.dina(n3254), .dinb(n3250), .dout(n3255));
  jand g2614(.dina(n3255), .dinb(n3235), .dout(n3256));
  jand g2615(.dina(n2628), .dinb(\in0[45] ), .dout(n3257));
  jand g2616(.dina(n2783), .dinb(\in1[45] ), .dout(n3258));
  jor  g2617(.dina(n3258), .dinb(n3257), .dout(n3259));
  jnot g2618(.din(n3259), .dout(n3260));
  jand g2619(.dina(n1556), .dinb(\in2[45] ), .dout(n3261));
  jand g2620(.dina(n1711), .dinb(\in3[45] ), .dout(n3262));
  jor  g2621(.dina(n3262), .dinb(n3261), .dout(n3263));
  jand g2622(.dina(n3263), .dinb(n3260), .dout(n3264));
  jand g2623(.dina(n2628), .dinb(\in0[47] ), .dout(n3265));
  jand g2624(.dina(n2783), .dinb(\in1[47] ), .dout(n3266));
  jor  g2625(.dina(n3266), .dinb(n3265), .dout(n3267));
  jnot g2626(.din(n3267), .dout(n3268));
  jand g2627(.dina(n1556), .dinb(\in2[47] ), .dout(n3269));
  jand g2628(.dina(n1711), .dinb(\in3[47] ), .dout(n3270));
  jor  g2629(.dina(n3270), .dinb(n3269), .dout(n3271));
  jand g2630(.dina(n3271), .dinb(n3268), .dout(n3272));
  jand g2631(.dina(n1556), .dinb(\in2[46] ), .dout(n3273));
  jand g2632(.dina(n1711), .dinb(\in3[46] ), .dout(n3274));
  jor  g2633(.dina(n3274), .dinb(n3273), .dout(n3275));
  jand g2634(.dina(n2628), .dinb(\in0[46] ), .dout(n3276));
  jand g2635(.dina(n2783), .dinb(\in1[46] ), .dout(n3277));
  jor  g2636(.dina(n3277), .dinb(n3276), .dout(n3278));
  jnot g2637(.din(n3278), .dout(n3279));
  jand g2638(.dina(n3279), .dinb(n3275), .dout(n3280));
  jor  g2639(.dina(n3280), .dinb(n3272), .dout(n3281));
  jor  g2640(.dina(n3281), .dinb(n3264), .dout(n3282));
  jand g2641(.dina(n2628), .dinb(\in0[43] ), .dout(n3283));
  jand g2642(.dina(n2783), .dinb(\in1[43] ), .dout(n3284));
  jor  g2643(.dina(n3284), .dinb(n3283), .dout(n3285));
  jnot g2644(.din(n3285), .dout(n3286));
  jand g2645(.dina(n1556), .dinb(\in2[43] ), .dout(n3287));
  jand g2646(.dina(n1711), .dinb(\in3[43] ), .dout(n3288));
  jor  g2647(.dina(n3288), .dinb(n3287), .dout(n3289));
  jand g2648(.dina(n3289), .dinb(n3286), .dout(n3290));
  jand g2649(.dina(n2628), .dinb(\in0[42] ), .dout(n3291));
  jand g2650(.dina(n2783), .dinb(\in1[42] ), .dout(n3292));
  jor  g2651(.dina(n3292), .dinb(n3291), .dout(n3293));
  jnot g2652(.din(n3293), .dout(n3294));
  jand g2653(.dina(n1556), .dinb(\in2[42] ), .dout(n3295));
  jand g2654(.dina(n1711), .dinb(\in3[42] ), .dout(n3296));
  jor  g2655(.dina(n3296), .dinb(n3295), .dout(n3297));
  jand g2656(.dina(n3297), .dinb(n3294), .dout(n3298));
  jor  g2657(.dina(n3298), .dinb(n3290), .dout(n3299));
  jand g2658(.dina(n2628), .dinb(\in0[44] ), .dout(n3300));
  jand g2659(.dina(n2783), .dinb(\in1[44] ), .dout(n3301));
  jor  g2660(.dina(n3301), .dinb(n3300), .dout(n3302));
  jnot g2661(.din(n3302), .dout(n3303));
  jand g2662(.dina(n1556), .dinb(\in2[44] ), .dout(n3304));
  jand g2663(.dina(n1711), .dinb(\in3[44] ), .dout(n3305));
  jor  g2664(.dina(n3305), .dinb(n3304), .dout(n3306));
  jand g2665(.dina(n3306), .dinb(n3303), .dout(n3307));
  jand g2666(.dina(n2628), .dinb(\in0[40] ), .dout(n3308));
  jand g2667(.dina(n2783), .dinb(\in1[40] ), .dout(n3309));
  jor  g2668(.dina(n3309), .dinb(n3308), .dout(n3310));
  jnot g2669(.din(n3310), .dout(n3311));
  jand g2670(.dina(n1556), .dinb(\in2[40] ), .dout(n3312));
  jand g2671(.dina(n1711), .dinb(\in3[40] ), .dout(n3313));
  jor  g2672(.dina(n3313), .dinb(n3312), .dout(n3314));
  jand g2673(.dina(n3314), .dinb(n3311), .dout(n3315));
  jand g2674(.dina(n2628), .dinb(\in0[41] ), .dout(n3316));
  jand g2675(.dina(n2783), .dinb(\in1[41] ), .dout(n3317));
  jor  g2676(.dina(n3317), .dinb(n3316), .dout(n3318));
  jnot g2677(.din(n3318), .dout(n3319));
  jand g2678(.dina(n1556), .dinb(\in2[41] ), .dout(n3320));
  jand g2679(.dina(n1711), .dinb(\in3[41] ), .dout(n3321));
  jor  g2680(.dina(n3321), .dinb(n3320), .dout(n3322));
  jand g2681(.dina(n3322), .dinb(n3319), .dout(n3323));
  jor  g2682(.dina(n3323), .dinb(n3315), .dout(n3324));
  jor  g2683(.dina(n3324), .dinb(n3307), .dout(n3325));
  jor  g2684(.dina(n3325), .dinb(n3299), .dout(n3326));
  jor  g2685(.dina(n3326), .dinb(n3282), .dout(n3327));
  jor  g2686(.dina(n3327), .dinb(n3256), .dout(n3328));
  jor  g2687(.dina(n3289), .dinb(n3286), .dout(n3329));
  jor  g2688(.dina(n3314), .dinb(n3311), .dout(n3330));
  jor  g2689(.dina(n3330), .dinb(n3323), .dout(n3331));
  jor  g2690(.dina(n3322), .dinb(n3319), .dout(n3332));
  jor  g2691(.dina(n3297), .dinb(n3294), .dout(n3333));
  jand g2692(.dina(n3333), .dinb(n3332), .dout(n3334));
  jand g2693(.dina(n3334), .dinb(n3331), .dout(n3335));
  jor  g2694(.dina(n3335), .dinb(n3299), .dout(n3336));
  jand g2695(.dina(n3336), .dinb(n3329), .dout(n3337));
  jor  g2696(.dina(n3337), .dinb(n3307), .dout(n3338));
  jor  g2697(.dina(n3306), .dinb(n3303), .dout(n3339));
  jor  g2698(.dina(n3263), .dinb(n3260), .dout(n3340));
  jand g2699(.dina(n3340), .dinb(n3339), .dout(n3341));
  jand g2700(.dina(n3341), .dinb(n3338), .dout(n3342));
  jor  g2701(.dina(n3342), .dinb(n3282), .dout(n3343));
  jor  g2702(.dina(n3279), .dinb(n3275), .dout(n3344));
  jor  g2703(.dina(n3344), .dinb(n3272), .dout(n3345));
  jor  g2704(.dina(n3271), .dinb(n3268), .dout(n3346));
  jand g2705(.dina(n3346), .dinb(n3345), .dout(n3347));
  jand g2706(.dina(n3347), .dinb(n3343), .dout(n3348));
  jand g2707(.dina(n3348), .dinb(n3328), .dout(n3349));
  jand g2708(.dina(n2628), .dinb(\in0[51] ), .dout(n3350));
  jand g2709(.dina(n2783), .dinb(\in1[51] ), .dout(n3351));
  jor  g2710(.dina(n3351), .dinb(n3350), .dout(n3352));
  jnot g2711(.din(n3352), .dout(n3353));
  jand g2712(.dina(n1556), .dinb(\in2[51] ), .dout(n3354));
  jand g2713(.dina(n1711), .dinb(\in3[51] ), .dout(n3355));
  jor  g2714(.dina(n3355), .dinb(n3354), .dout(n3356));
  jand g2715(.dina(n3356), .dinb(n3353), .dout(n3357));
  jand g2716(.dina(n2628), .dinb(\in0[49] ), .dout(n3358));
  jand g2717(.dina(n2783), .dinb(\in1[49] ), .dout(n3359));
  jor  g2718(.dina(n3359), .dinb(n3358), .dout(n3360));
  jnot g2719(.din(n3360), .dout(n3361));
  jand g2720(.dina(n1556), .dinb(\in2[49] ), .dout(n3362));
  jand g2721(.dina(n1711), .dinb(\in3[49] ), .dout(n3363));
  jor  g2722(.dina(n3363), .dinb(n3362), .dout(n3364));
  jand g2723(.dina(n3364), .dinb(n3361), .dout(n3365));
  jand g2724(.dina(n1556), .dinb(\in2[50] ), .dout(n3366));
  jand g2725(.dina(n1711), .dinb(\in3[50] ), .dout(n3367));
  jor  g2726(.dina(n3367), .dinb(n3366), .dout(n3368));
  jand g2727(.dina(n2628), .dinb(\in0[50] ), .dout(n3369));
  jand g2728(.dina(n2783), .dinb(\in1[50] ), .dout(n3370));
  jor  g2729(.dina(n3370), .dinb(n3369), .dout(n3371));
  jnot g2730(.din(n3371), .dout(n3372));
  jand g2731(.dina(n3372), .dinb(n3368), .dout(n3373));
  jor  g2732(.dina(n3373), .dinb(n3365), .dout(n3374));
  jor  g2733(.dina(n3374), .dinb(n3357), .dout(n3375));
  jand g2734(.dina(n2628), .dinb(\in0[53] ), .dout(n3376));
  jand g2735(.dina(n2783), .dinb(\in1[53] ), .dout(n3377));
  jor  g2736(.dina(n3377), .dinb(n3376), .dout(n3378));
  jnot g2737(.din(n3378), .dout(n3379));
  jand g2738(.dina(n1556), .dinb(\in2[53] ), .dout(n3380));
  jand g2739(.dina(n1711), .dinb(\in3[53] ), .dout(n3381));
  jor  g2740(.dina(n3381), .dinb(n3380), .dout(n3382));
  jand g2741(.dina(n3382), .dinb(n3379), .dout(n3383));
  jnot g2742(.din(n3383), .dout(n3384));
  jand g2743(.dina(n2628), .dinb(\in0[52] ), .dout(n3385));
  jand g2744(.dina(n2783), .dinb(\in1[52] ), .dout(n3386));
  jor  g2745(.dina(n3386), .dinb(n3385), .dout(n3387));
  jand g2746(.dina(n3387), .dinb(n3384), .dout(n3388));
  jand g2747(.dina(n1556), .dinb(\in2[52] ), .dout(n3389));
  jand g2748(.dina(n1711), .dinb(\in3[52] ), .dout(n3390));
  jor  g2749(.dina(n3390), .dinb(n3389), .dout(n3391));
  jnot g2750(.din(n3391), .dout(n3392));
  jand g2751(.dina(n3392), .dinb(n3384), .dout(n3393));
  jor  g2752(.dina(n3393), .dinb(n3388), .dout(n3394));
  jnot g2753(.din(n3394), .dout(n3395));
  jand g2754(.dina(n2628), .dinb(\in0[55] ), .dout(n3396));
  jand g2755(.dina(n2783), .dinb(\in1[55] ), .dout(n3397));
  jor  g2756(.dina(n3397), .dinb(n3396), .dout(n3398));
  jnot g2757(.din(n3398), .dout(n3399));
  jand g2758(.dina(n1556), .dinb(\in2[55] ), .dout(n3400));
  jand g2759(.dina(n1711), .dinb(\in3[55] ), .dout(n3401));
  jor  g2760(.dina(n3401), .dinb(n3400), .dout(n3402));
  jand g2761(.dina(n3402), .dinb(n3399), .dout(n3403));
  jand g2762(.dina(n1556), .dinb(\in2[54] ), .dout(n3404));
  jand g2763(.dina(n1711), .dinb(\in3[54] ), .dout(n3405));
  jor  g2764(.dina(n3405), .dinb(n3404), .dout(n3406));
  jand g2765(.dina(n2628), .dinb(\in0[54] ), .dout(n3407));
  jand g2766(.dina(n2783), .dinb(\in1[54] ), .dout(n3408));
  jor  g2767(.dina(n3408), .dinb(n3407), .dout(n3409));
  jnot g2768(.din(n3409), .dout(n3410));
  jand g2769(.dina(n3410), .dinb(n3406), .dout(n3411));
  jor  g2770(.dina(n3411), .dinb(n3403), .dout(n3412));
  jand g2771(.dina(n1556), .dinb(\in2[48] ), .dout(n3413));
  jand g2772(.dina(n1711), .dinb(\in3[48] ), .dout(n3414));
  jor  g2773(.dina(n3414), .dinb(n3413), .dout(n3415));
  jand g2774(.dina(n2628), .dinb(\in0[48] ), .dout(n3416));
  jand g2775(.dina(n2783), .dinb(\in1[48] ), .dout(n3417));
  jor  g2776(.dina(n3417), .dinb(n3416), .dout(n3418));
  jnot g2777(.din(n3418), .dout(n3419));
  jand g2778(.dina(n3419), .dinb(n3415), .dout(n3420));
  jor  g2779(.dina(n3420), .dinb(n3412), .dout(n3421));
  jor  g2780(.dina(n3421), .dinb(n3395), .dout(n3422));
  jor  g2781(.dina(n3422), .dinb(n3375), .dout(n3423));
  jor  g2782(.dina(n3423), .dinb(n3349), .dout(n3424));
  jor  g2783(.dina(n3402), .dinb(n3399), .dout(n3425));
  jor  g2784(.dina(n3419), .dinb(n3415), .dout(n3426));
  jor  g2785(.dina(n3364), .dinb(n3361), .dout(n3427));
  jand g2786(.dina(n3427), .dinb(n3426), .dout(n3428));
  jor  g2787(.dina(n3428), .dinb(n3375), .dout(n3429));
  jor  g2788(.dina(n3372), .dinb(n3368), .dout(n3430));
  jor  g2789(.dina(n3430), .dinb(n3357), .dout(n3431));
  jor  g2790(.dina(n3356), .dinb(n3353), .dout(n3432));
  jand g2791(.dina(n3432), .dinb(n3431), .dout(n3433));
  jand g2792(.dina(n3433), .dinb(n3429), .dout(n3434));
  jor  g2793(.dina(n3434), .dinb(n3395), .dout(n3435));
  jand g2794(.dina(n3392), .dinb(n3388), .dout(n3436));
  jnot g2795(.din(n3436), .dout(n3437));
  jor  g2796(.dina(n3382), .dinb(n3379), .dout(n3438));
  jor  g2797(.dina(n3410), .dinb(n3406), .dout(n3439));
  jand g2798(.dina(n3439), .dinb(n3438), .dout(n3440));
  jand g2799(.dina(n3440), .dinb(n3437), .dout(n3441));
  jand g2800(.dina(n3441), .dinb(n3435), .dout(n3442));
  jor  g2801(.dina(n3442), .dinb(n3412), .dout(n3443));
  jand g2802(.dina(n3443), .dinb(n3425), .dout(n3444));
  jand g2803(.dina(n3444), .dinb(n3424), .dout(n3445));
  jand g2804(.dina(n2628), .dinb(\in0[61] ), .dout(n3446));
  jand g2805(.dina(n2783), .dinb(\in1[61] ), .dout(n3447));
  jor  g2806(.dina(n3447), .dinb(n3446), .dout(n3448));
  jnot g2807(.din(n3448), .dout(n3449));
  jand g2808(.dina(n1556), .dinb(\in2[61] ), .dout(n3450));
  jand g2809(.dina(n1711), .dinb(\in3[61] ), .dout(n3451));
  jor  g2810(.dina(n3451), .dinb(n3450), .dout(n3452));
  jand g2811(.dina(n3452), .dinb(n3449), .dout(n3453));
  jand g2812(.dina(n2628), .dinb(\in0[63] ), .dout(n3454));
  jand g2813(.dina(n2783), .dinb(\in1[63] ), .dout(n3455));
  jor  g2814(.dina(n3455), .dinb(n3454), .dout(n3456));
  jnot g2815(.din(n3456), .dout(n3457));
  jand g2816(.dina(n1556), .dinb(\in2[63] ), .dout(n3458));
  jand g2817(.dina(n1711), .dinb(\in3[63] ), .dout(n3459));
  jor  g2818(.dina(n3459), .dinb(n3458), .dout(n3460));
  jand g2819(.dina(n3460), .dinb(n3457), .dout(n3461));
  jand g2820(.dina(n1556), .dinb(\in2[62] ), .dout(n3462));
  jand g2821(.dina(n1711), .dinb(\in3[62] ), .dout(n3463));
  jor  g2822(.dina(n3463), .dinb(n3462), .dout(n3464));
  jand g2823(.dina(n2628), .dinb(\in0[62] ), .dout(n3465));
  jand g2824(.dina(n2783), .dinb(\in1[62] ), .dout(n3466));
  jor  g2825(.dina(n3466), .dinb(n3465), .dout(n3467));
  jnot g2826(.din(n3467), .dout(n3468));
  jand g2827(.dina(n3468), .dinb(n3464), .dout(n3469));
  jor  g2828(.dina(n3469), .dinb(n3461), .dout(n3470));
  jor  g2829(.dina(n3470), .dinb(n3453), .dout(n3471));
  jand g2830(.dina(n2628), .dinb(\in0[59] ), .dout(n3472));
  jand g2831(.dina(n2783), .dinb(\in1[59] ), .dout(n3473));
  jor  g2832(.dina(n3473), .dinb(n3472), .dout(n3474));
  jnot g2833(.din(n3474), .dout(n3475));
  jand g2834(.dina(n1556), .dinb(\in2[59] ), .dout(n3476));
  jand g2835(.dina(n1711), .dinb(\in3[59] ), .dout(n3477));
  jor  g2836(.dina(n3477), .dinb(n3476), .dout(n3478));
  jand g2837(.dina(n3478), .dinb(n3475), .dout(n3479));
  jand g2838(.dina(n2628), .dinb(\in0[58] ), .dout(n3480));
  jand g2839(.dina(n2783), .dinb(\in1[58] ), .dout(n3481));
  jor  g2840(.dina(n3481), .dinb(n3480), .dout(n3482));
  jnot g2841(.din(n3482), .dout(n3483));
  jand g2842(.dina(n1556), .dinb(\in2[58] ), .dout(n3484));
  jand g2843(.dina(n1711), .dinb(\in3[58] ), .dout(n3485));
  jor  g2844(.dina(n3485), .dinb(n3484), .dout(n3486));
  jand g2845(.dina(n3486), .dinb(n3483), .dout(n3487));
  jor  g2846(.dina(n3487), .dinb(n3479), .dout(n3488));
  jand g2847(.dina(n2628), .dinb(\in0[60] ), .dout(n3489));
  jand g2848(.dina(n2783), .dinb(\in1[60] ), .dout(n3490));
  jor  g2849(.dina(n3490), .dinb(n3489), .dout(n3491));
  jnot g2850(.din(n3491), .dout(n3492));
  jand g2851(.dina(n1556), .dinb(\in2[60] ), .dout(n3493));
  jand g2852(.dina(n1711), .dinb(\in3[60] ), .dout(n3494));
  jor  g2853(.dina(n3494), .dinb(n3493), .dout(n3495));
  jand g2854(.dina(n3495), .dinb(n3492), .dout(n3496));
  jand g2855(.dina(n2628), .dinb(\in0[56] ), .dout(n3497));
  jand g2856(.dina(n2783), .dinb(\in1[56] ), .dout(n3498));
  jor  g2857(.dina(n3498), .dinb(n3497), .dout(n3499));
  jnot g2858(.din(n3499), .dout(n3500));
  jand g2859(.dina(n1556), .dinb(\in2[56] ), .dout(n3501));
  jand g2860(.dina(n1711), .dinb(\in3[56] ), .dout(n3502));
  jor  g2861(.dina(n3502), .dinb(n3501), .dout(n3503));
  jand g2862(.dina(n3503), .dinb(n3500), .dout(n3504));
  jand g2863(.dina(n2628), .dinb(\in0[57] ), .dout(n3505));
  jand g2864(.dina(n2783), .dinb(\in1[57] ), .dout(n3506));
  jor  g2865(.dina(n3506), .dinb(n3505), .dout(n3507));
  jnot g2866(.din(n3507), .dout(n3508));
  jand g2867(.dina(n1556), .dinb(\in2[57] ), .dout(n3509));
  jand g2868(.dina(n1711), .dinb(\in3[57] ), .dout(n3510));
  jor  g2869(.dina(n3510), .dinb(n3509), .dout(n3511));
  jand g2870(.dina(n3511), .dinb(n3508), .dout(n3512));
  jor  g2871(.dina(n3512), .dinb(n3504), .dout(n3513));
  jor  g2872(.dina(n3513), .dinb(n3496), .dout(n3514));
  jor  g2873(.dina(n3514), .dinb(n3488), .dout(n3515));
  jor  g2874(.dina(n3515), .dinb(n3471), .dout(n3516));
  jor  g2875(.dina(n3516), .dinb(n3445), .dout(n3517));
  jor  g2876(.dina(n3478), .dinb(n3475), .dout(n3518));
  jor  g2877(.dina(n3503), .dinb(n3500), .dout(n3519));
  jor  g2878(.dina(n3519), .dinb(n3512), .dout(n3520));
  jor  g2879(.dina(n3511), .dinb(n3508), .dout(n3521));
  jor  g2880(.dina(n3486), .dinb(n3483), .dout(n3522));
  jand g2881(.dina(n3522), .dinb(n3521), .dout(n3523));
  jand g2882(.dina(n3523), .dinb(n3520), .dout(n3524));
  jor  g2883(.dina(n3524), .dinb(n3488), .dout(n3525));
  jand g2884(.dina(n3525), .dinb(n3518), .dout(n3526));
  jor  g2885(.dina(n3526), .dinb(n3496), .dout(n3527));
  jor  g2886(.dina(n3495), .dinb(n3492), .dout(n3528));
  jor  g2887(.dina(n3452), .dinb(n3449), .dout(n3529));
  jand g2888(.dina(n3529), .dinb(n3528), .dout(n3530));
  jand g2889(.dina(n3530), .dinb(n3527), .dout(n3531));
  jor  g2890(.dina(n3531), .dinb(n3471), .dout(n3532));
  jor  g2891(.dina(n3468), .dinb(n3464), .dout(n3533));
  jor  g2892(.dina(n3533), .dinb(n3461), .dout(n3534));
  jor  g2893(.dina(n3460), .dinb(n3457), .dout(n3535));
  jand g2894(.dina(n3535), .dinb(n3534), .dout(n3536));
  jand g2895(.dina(n3536), .dinb(n3532), .dout(n3537));
  jand g2896(.dina(n3537), .dinb(n3517), .dout(n3538));
  jand g2897(.dina(n2628), .dinb(\in0[67] ), .dout(n3539));
  jand g2898(.dina(n2783), .dinb(\in1[67] ), .dout(n3540));
  jor  g2899(.dina(n3540), .dinb(n3539), .dout(n3541));
  jnot g2900(.din(n3541), .dout(n3542));
  jand g2901(.dina(n1556), .dinb(\in2[67] ), .dout(n3543));
  jand g2902(.dina(n1711), .dinb(\in3[67] ), .dout(n3544));
  jor  g2903(.dina(n3544), .dinb(n3543), .dout(n3545));
  jand g2904(.dina(n3545), .dinb(n3542), .dout(n3546));
  jand g2905(.dina(n1556), .dinb(\in2[66] ), .dout(n3547));
  jand g2906(.dina(n1711), .dinb(\in3[66] ), .dout(n3548));
  jor  g2907(.dina(n3548), .dinb(n3547), .dout(n3549));
  jand g2908(.dina(n2628), .dinb(\in0[66] ), .dout(n3550));
  jand g2909(.dina(n2783), .dinb(\in1[66] ), .dout(n3551));
  jor  g2910(.dina(n3551), .dinb(n3550), .dout(n3552));
  jnot g2911(.din(n3552), .dout(n3553));
  jand g2912(.dina(n3553), .dinb(n3549), .dout(n3554));
  jor  g2913(.dina(n3554), .dinb(n3546), .dout(n3555));
  jand g2914(.dina(n2628), .dinb(\in0[65] ), .dout(n3556));
  jand g2915(.dina(n2783), .dinb(\in1[65] ), .dout(n3557));
  jor  g2916(.dina(n3557), .dinb(n3556), .dout(n3558));
  jnot g2917(.din(n3558), .dout(n3559));
  jand g2918(.dina(n1556), .dinb(\in2[65] ), .dout(n3560));
  jand g2919(.dina(n1711), .dinb(\in3[65] ), .dout(n3561));
  jor  g2920(.dina(n3561), .dinb(n3560), .dout(n3562));
  jand g2921(.dina(n3562), .dinb(n3559), .dout(n3563));
  jand g2922(.dina(n1556), .dinb(\in2[64] ), .dout(n3564));
  jand g2923(.dina(n1711), .dinb(\in3[64] ), .dout(n3565));
  jor  g2924(.dina(n3565), .dinb(n3564), .dout(n3566));
  jand g2925(.dina(n2628), .dinb(\in0[64] ), .dout(n3567));
  jand g2926(.dina(n2783), .dinb(\in1[64] ), .dout(n3568));
  jor  g2927(.dina(n3568), .dinb(n3567), .dout(n3569));
  jnot g2928(.din(n3569), .dout(n3570));
  jand g2929(.dina(n3570), .dinb(n3566), .dout(n3571));
  jor  g2930(.dina(n3571), .dinb(n3563), .dout(n3572));
  jor  g2931(.dina(n3572), .dinb(n3555), .dout(n3573));
  jor  g2932(.dina(n3573), .dinb(n3538), .dout(n3574));
  jor  g2933(.dina(n3545), .dinb(n3542), .dout(n3575));
  jor  g2934(.dina(n3570), .dinb(n3566), .dout(n3576));
  jor  g2935(.dina(n3576), .dinb(n3563), .dout(n3577));
  jor  g2936(.dina(n3562), .dinb(n3559), .dout(n3578));
  jor  g2937(.dina(n3553), .dinb(n3549), .dout(n3579));
  jand g2938(.dina(n3579), .dinb(n3578), .dout(n3580));
  jand g2939(.dina(n3580), .dinb(n3577), .dout(n3581));
  jor  g2940(.dina(n3581), .dinb(n3555), .dout(n3582));
  jand g2941(.dina(n3582), .dinb(n3575), .dout(n3583));
  jand g2942(.dina(n3583), .dinb(n3574), .dout(n3584));
  jand g2943(.dina(n2628), .dinb(\in0[68] ), .dout(n3585));
  jand g2944(.dina(n2783), .dinb(\in1[68] ), .dout(n3586));
  jor  g2945(.dina(n3586), .dinb(n3585), .dout(n3587));
  jnot g2946(.din(n3587), .dout(n3588));
  jand g2947(.dina(n1556), .dinb(\in2[68] ), .dout(n3589));
  jand g2948(.dina(n1711), .dinb(\in3[68] ), .dout(n3590));
  jor  g2949(.dina(n3590), .dinb(n3589), .dout(n3591));
  jand g2950(.dina(n3591), .dinb(n3588), .dout(n3592));
  jand g2951(.dina(n2628), .dinb(\in0[69] ), .dout(n3593));
  jand g2952(.dina(n2783), .dinb(\in1[69] ), .dout(n3594));
  jor  g2953(.dina(n3594), .dinb(n3593), .dout(n3595));
  jnot g2954(.din(n3595), .dout(n3596));
  jand g2955(.dina(n1556), .dinb(\in2[69] ), .dout(n3597));
  jand g2956(.dina(n1711), .dinb(\in3[69] ), .dout(n3598));
  jor  g2957(.dina(n3598), .dinb(n3597), .dout(n3599));
  jand g2958(.dina(n3599), .dinb(n3596), .dout(n3600));
  jand g2959(.dina(n2628), .dinb(\in0[71] ), .dout(n3601));
  jand g2960(.dina(n2783), .dinb(\in1[71] ), .dout(n3602));
  jor  g2961(.dina(n3602), .dinb(n3601), .dout(n3603));
  jnot g2962(.din(n3603), .dout(n3604));
  jand g2963(.dina(n1556), .dinb(\in2[71] ), .dout(n3605));
  jand g2964(.dina(n1711), .dinb(\in3[71] ), .dout(n3606));
  jor  g2965(.dina(n3606), .dinb(n3605), .dout(n3607));
  jand g2966(.dina(n3607), .dinb(n3604), .dout(n3608));
  jand g2967(.dina(n1556), .dinb(\in2[70] ), .dout(n3609));
  jand g2968(.dina(n1711), .dinb(\in3[70] ), .dout(n3610));
  jor  g2969(.dina(n3610), .dinb(n3609), .dout(n3611));
  jand g2970(.dina(n2628), .dinb(\in0[70] ), .dout(n3612));
  jand g2971(.dina(n2783), .dinb(\in1[70] ), .dout(n3613));
  jor  g2972(.dina(n3613), .dinb(n3612), .dout(n3614));
  jnot g2973(.din(n3614), .dout(n3615));
  jand g2974(.dina(n3615), .dinb(n3611), .dout(n3616));
  jor  g2975(.dina(n3616), .dinb(n3608), .dout(n3617));
  jor  g2976(.dina(n3617), .dinb(n3600), .dout(n3618));
  jor  g2977(.dina(n3618), .dinb(n3592), .dout(n3619));
  jor  g2978(.dina(n3619), .dinb(n3584), .dout(n3620));
  jor  g2979(.dina(n3599), .dinb(n3596), .dout(n3621));
  jor  g2980(.dina(n3591), .dinb(n3588), .dout(n3622));
  jand g2981(.dina(n3622), .dinb(n3621), .dout(n3623));
  jor  g2982(.dina(n3623), .dinb(n3618), .dout(n3624));
  jor  g2983(.dina(n3607), .dinb(n3604), .dout(n3625));
  jor  g2984(.dina(n3615), .dinb(n3611), .dout(n3626));
  jor  g2985(.dina(n3626), .dinb(n3608), .dout(n3627));
  jand g2986(.dina(n3627), .dinb(n3625), .dout(n3628));
  jand g2987(.dina(n3628), .dinb(n3624), .dout(n3629));
  jand g2988(.dina(n3629), .dinb(n3620), .dout(n3630));
  jand g2989(.dina(n2628), .dinb(\in0[75] ), .dout(n3631));
  jand g2990(.dina(n2783), .dinb(\in1[75] ), .dout(n3632));
  jor  g2991(.dina(n3632), .dinb(n3631), .dout(n3633));
  jnot g2992(.din(n3633), .dout(n3634));
  jand g2993(.dina(n1556), .dinb(\in2[75] ), .dout(n3635));
  jand g2994(.dina(n1711), .dinb(\in3[75] ), .dout(n3636));
  jor  g2995(.dina(n3636), .dinb(n3635), .dout(n3637));
  jand g2996(.dina(n3637), .dinb(n3634), .dout(n3638));
  jand g2997(.dina(n1556), .dinb(\in2[74] ), .dout(n3639));
  jand g2998(.dina(n1711), .dinb(\in3[74] ), .dout(n3640));
  jor  g2999(.dina(n3640), .dinb(n3639), .dout(n3641));
  jand g3000(.dina(n2628), .dinb(\in0[74] ), .dout(n3642));
  jand g3001(.dina(n2783), .dinb(\in1[74] ), .dout(n3643));
  jor  g3002(.dina(n3643), .dinb(n3642), .dout(n3644));
  jnot g3003(.din(n3644), .dout(n3645));
  jand g3004(.dina(n3645), .dinb(n3641), .dout(n3646));
  jor  g3005(.dina(n3646), .dinb(n3638), .dout(n3647));
  jand g3006(.dina(n2628), .dinb(\in0[73] ), .dout(n3648));
  jand g3007(.dina(n2783), .dinb(\in1[73] ), .dout(n3649));
  jor  g3008(.dina(n3649), .dinb(n3648), .dout(n3650));
  jnot g3009(.din(n3650), .dout(n3651));
  jand g3010(.dina(n1556), .dinb(\in2[73] ), .dout(n3652));
  jand g3011(.dina(n1711), .dinb(\in3[73] ), .dout(n3653));
  jor  g3012(.dina(n3653), .dinb(n3652), .dout(n3654));
  jand g3013(.dina(n3654), .dinb(n3651), .dout(n3655));
  jand g3014(.dina(n1556), .dinb(\in2[72] ), .dout(n3656));
  jand g3015(.dina(n1711), .dinb(\in3[72] ), .dout(n3657));
  jor  g3016(.dina(n3657), .dinb(n3656), .dout(n3658));
  jand g3017(.dina(n2628), .dinb(\in0[72] ), .dout(n3659));
  jand g3018(.dina(n2783), .dinb(\in1[72] ), .dout(n3660));
  jor  g3019(.dina(n3660), .dinb(n3659), .dout(n3661));
  jnot g3020(.din(n3661), .dout(n3662));
  jand g3021(.dina(n3662), .dinb(n3658), .dout(n3663));
  jor  g3022(.dina(n3663), .dinb(n3655), .dout(n3664));
  jor  g3023(.dina(n3664), .dinb(n3647), .dout(n3665));
  jor  g3024(.dina(n3665), .dinb(n3630), .dout(n3666));
  jor  g3025(.dina(n3637), .dinb(n3634), .dout(n3667));
  jor  g3026(.dina(n3662), .dinb(n3658), .dout(n3668));
  jor  g3027(.dina(n3668), .dinb(n3655), .dout(n3669));
  jor  g3028(.dina(n3654), .dinb(n3651), .dout(n3670));
  jor  g3029(.dina(n3645), .dinb(n3641), .dout(n3671));
  jand g3030(.dina(n3671), .dinb(n3670), .dout(n3672));
  jand g3031(.dina(n3672), .dinb(n3669), .dout(n3673));
  jor  g3032(.dina(n3673), .dinb(n3647), .dout(n3674));
  jand g3033(.dina(n3674), .dinb(n3667), .dout(n3675));
  jand g3034(.dina(n3675), .dinb(n3666), .dout(n3676));
  jand g3035(.dina(n2628), .dinb(\in0[76] ), .dout(n3677));
  jand g3036(.dina(n2783), .dinb(\in1[76] ), .dout(n3678));
  jor  g3037(.dina(n3678), .dinb(n3677), .dout(n3679));
  jnot g3038(.din(n3679), .dout(n3680));
  jand g3039(.dina(n1556), .dinb(\in2[76] ), .dout(n3681));
  jand g3040(.dina(n1711), .dinb(\in3[76] ), .dout(n3682));
  jor  g3041(.dina(n3682), .dinb(n3681), .dout(n3683));
  jand g3042(.dina(n3683), .dinb(n3680), .dout(n3684));
  jand g3043(.dina(n2628), .dinb(\in0[77] ), .dout(n3685));
  jand g3044(.dina(n2783), .dinb(\in1[77] ), .dout(n3686));
  jor  g3045(.dina(n3686), .dinb(n3685), .dout(n3687));
  jnot g3046(.din(n3687), .dout(n3688));
  jand g3047(.dina(n1556), .dinb(\in2[77] ), .dout(n3689));
  jand g3048(.dina(n1711), .dinb(\in3[77] ), .dout(n3690));
  jor  g3049(.dina(n3690), .dinb(n3689), .dout(n3691));
  jand g3050(.dina(n3691), .dinb(n3688), .dout(n3692));
  jand g3051(.dina(n2628), .dinb(\in0[79] ), .dout(n3693));
  jand g3052(.dina(n2783), .dinb(\in1[79] ), .dout(n3694));
  jor  g3053(.dina(n3694), .dinb(n3693), .dout(n3695));
  jnot g3054(.din(n3695), .dout(n3696));
  jand g3055(.dina(n1556), .dinb(\in2[79] ), .dout(n3697));
  jand g3056(.dina(n1711), .dinb(\in3[79] ), .dout(n3698));
  jor  g3057(.dina(n3698), .dinb(n3697), .dout(n3699));
  jand g3058(.dina(n3699), .dinb(n3696), .dout(n3700));
  jand g3059(.dina(n1556), .dinb(\in2[78] ), .dout(n3701));
  jand g3060(.dina(n1711), .dinb(\in3[78] ), .dout(n3702));
  jor  g3061(.dina(n3702), .dinb(n3701), .dout(n3703));
  jand g3062(.dina(n2628), .dinb(\in0[78] ), .dout(n3704));
  jand g3063(.dina(n2783), .dinb(\in1[78] ), .dout(n3705));
  jor  g3064(.dina(n3705), .dinb(n3704), .dout(n3706));
  jnot g3065(.din(n3706), .dout(n3707));
  jand g3066(.dina(n3707), .dinb(n3703), .dout(n3708));
  jor  g3067(.dina(n3708), .dinb(n3700), .dout(n3709));
  jor  g3068(.dina(n3709), .dinb(n3692), .dout(n3710));
  jor  g3069(.dina(n3710), .dinb(n3684), .dout(n3711));
  jor  g3070(.dina(n3711), .dinb(n3676), .dout(n3712));
  jor  g3071(.dina(n3691), .dinb(n3688), .dout(n3713));
  jor  g3072(.dina(n3683), .dinb(n3680), .dout(n3714));
  jand g3073(.dina(n3714), .dinb(n3713), .dout(n3715));
  jor  g3074(.dina(n3715), .dinb(n3710), .dout(n3716));
  jor  g3075(.dina(n3699), .dinb(n3696), .dout(n3717));
  jor  g3076(.dina(n3707), .dinb(n3703), .dout(n3718));
  jor  g3077(.dina(n3718), .dinb(n3700), .dout(n3719));
  jand g3078(.dina(n3719), .dinb(n3717), .dout(n3720));
  jand g3079(.dina(n3720), .dinb(n3716), .dout(n3721));
  jand g3080(.dina(n3721), .dinb(n3712), .dout(n3722));
  jand g3081(.dina(n2628), .dinb(\in0[83] ), .dout(n3723));
  jand g3082(.dina(n2783), .dinb(\in1[83] ), .dout(n3724));
  jor  g3083(.dina(n3724), .dinb(n3723), .dout(n3725));
  jnot g3084(.din(n3725), .dout(n3726));
  jand g3085(.dina(n1556), .dinb(\in2[83] ), .dout(n3727));
  jand g3086(.dina(n1711), .dinb(\in3[83] ), .dout(n3728));
  jor  g3087(.dina(n3728), .dinb(n3727), .dout(n3729));
  jand g3088(.dina(n3729), .dinb(n3726), .dout(n3730));
  jand g3089(.dina(n1556), .dinb(\in2[82] ), .dout(n3731));
  jand g3090(.dina(n1711), .dinb(\in3[82] ), .dout(n3732));
  jor  g3091(.dina(n3732), .dinb(n3731), .dout(n3733));
  jand g3092(.dina(n2628), .dinb(\in0[82] ), .dout(n3734));
  jand g3093(.dina(n2783), .dinb(\in1[82] ), .dout(n3735));
  jor  g3094(.dina(n3735), .dinb(n3734), .dout(n3736));
  jnot g3095(.din(n3736), .dout(n3737));
  jand g3096(.dina(n3737), .dinb(n3733), .dout(n3738));
  jor  g3097(.dina(n3738), .dinb(n3730), .dout(n3739));
  jand g3098(.dina(n2628), .dinb(\in0[81] ), .dout(n3740));
  jand g3099(.dina(n2783), .dinb(\in1[81] ), .dout(n3741));
  jor  g3100(.dina(n3741), .dinb(n3740), .dout(n3742));
  jnot g3101(.din(n3742), .dout(n3743));
  jand g3102(.dina(n1556), .dinb(\in2[81] ), .dout(n3744));
  jand g3103(.dina(n1711), .dinb(\in3[81] ), .dout(n3745));
  jor  g3104(.dina(n3745), .dinb(n3744), .dout(n3746));
  jand g3105(.dina(n3746), .dinb(n3743), .dout(n3747));
  jand g3106(.dina(n1556), .dinb(\in2[80] ), .dout(n3748));
  jand g3107(.dina(n1711), .dinb(\in3[80] ), .dout(n3749));
  jor  g3108(.dina(n3749), .dinb(n3748), .dout(n3750));
  jand g3109(.dina(n2628), .dinb(\in0[80] ), .dout(n3751));
  jand g3110(.dina(n2783), .dinb(\in1[80] ), .dout(n3752));
  jor  g3111(.dina(n3752), .dinb(n3751), .dout(n3753));
  jnot g3112(.din(n3753), .dout(n3754));
  jand g3113(.dina(n3754), .dinb(n3750), .dout(n3755));
  jor  g3114(.dina(n3755), .dinb(n3747), .dout(n3756));
  jor  g3115(.dina(n3756), .dinb(n3739), .dout(n3757));
  jor  g3116(.dina(n3757), .dinb(n3722), .dout(n3758));
  jor  g3117(.dina(n3729), .dinb(n3726), .dout(n3759));
  jor  g3118(.dina(n3754), .dinb(n3750), .dout(n3760));
  jor  g3119(.dina(n3760), .dinb(n3747), .dout(n3761));
  jor  g3120(.dina(n3746), .dinb(n3743), .dout(n3762));
  jor  g3121(.dina(n3737), .dinb(n3733), .dout(n3763));
  jand g3122(.dina(n3763), .dinb(n3762), .dout(n3764));
  jand g3123(.dina(n3764), .dinb(n3761), .dout(n3765));
  jor  g3124(.dina(n3765), .dinb(n3739), .dout(n3766));
  jand g3125(.dina(n3766), .dinb(n3759), .dout(n3767));
  jand g3126(.dina(n3767), .dinb(n3758), .dout(n3768));
  jand g3127(.dina(n2628), .dinb(\in0[84] ), .dout(n3769));
  jand g3128(.dina(n2783), .dinb(\in1[84] ), .dout(n3770));
  jor  g3129(.dina(n3770), .dinb(n3769), .dout(n3771));
  jnot g3130(.din(n3771), .dout(n3772));
  jand g3131(.dina(n1556), .dinb(\in2[84] ), .dout(n3773));
  jand g3132(.dina(n1711), .dinb(\in3[84] ), .dout(n3774));
  jor  g3133(.dina(n3774), .dinb(n3773), .dout(n3775));
  jand g3134(.dina(n3775), .dinb(n3772), .dout(n3776));
  jand g3135(.dina(n2628), .dinb(\in0[85] ), .dout(n3777));
  jand g3136(.dina(n2783), .dinb(\in1[85] ), .dout(n3778));
  jor  g3137(.dina(n3778), .dinb(n3777), .dout(n3779));
  jnot g3138(.din(n3779), .dout(n3780));
  jand g3139(.dina(n1556), .dinb(\in2[85] ), .dout(n3781));
  jand g3140(.dina(n1711), .dinb(\in3[85] ), .dout(n3782));
  jor  g3141(.dina(n3782), .dinb(n3781), .dout(n3783));
  jand g3142(.dina(n3783), .dinb(n3780), .dout(n3784));
  jand g3143(.dina(n2628), .dinb(\in0[87] ), .dout(n3785));
  jand g3144(.dina(n2783), .dinb(\in1[87] ), .dout(n3786));
  jor  g3145(.dina(n3786), .dinb(n3785), .dout(n3787));
  jnot g3146(.din(n3787), .dout(n3788));
  jand g3147(.dina(n1556), .dinb(\in2[87] ), .dout(n3789));
  jand g3148(.dina(n1711), .dinb(\in3[87] ), .dout(n3790));
  jor  g3149(.dina(n3790), .dinb(n3789), .dout(n3791));
  jand g3150(.dina(n3791), .dinb(n3788), .dout(n3792));
  jand g3151(.dina(n1556), .dinb(\in2[86] ), .dout(n3793));
  jand g3152(.dina(n1711), .dinb(\in3[86] ), .dout(n3794));
  jor  g3153(.dina(n3794), .dinb(n3793), .dout(n3795));
  jand g3154(.dina(n2628), .dinb(\in0[86] ), .dout(n3796));
  jand g3155(.dina(n2783), .dinb(\in1[86] ), .dout(n3797));
  jor  g3156(.dina(n3797), .dinb(n3796), .dout(n3798));
  jnot g3157(.din(n3798), .dout(n3799));
  jand g3158(.dina(n3799), .dinb(n3795), .dout(n3800));
  jor  g3159(.dina(n3800), .dinb(n3792), .dout(n3801));
  jor  g3160(.dina(n3801), .dinb(n3784), .dout(n3802));
  jor  g3161(.dina(n3802), .dinb(n3776), .dout(n3803));
  jor  g3162(.dina(n3803), .dinb(n3768), .dout(n3804));
  jor  g3163(.dina(n3783), .dinb(n3780), .dout(n3805));
  jor  g3164(.dina(n3775), .dinb(n3772), .dout(n3806));
  jand g3165(.dina(n3806), .dinb(n3805), .dout(n3807));
  jor  g3166(.dina(n3807), .dinb(n3802), .dout(n3808));
  jor  g3167(.dina(n3791), .dinb(n3788), .dout(n3809));
  jor  g3168(.dina(n3799), .dinb(n3795), .dout(n3810));
  jor  g3169(.dina(n3810), .dinb(n3792), .dout(n3811));
  jand g3170(.dina(n3811), .dinb(n3809), .dout(n3812));
  jand g3171(.dina(n3812), .dinb(n3808), .dout(n3813));
  jand g3172(.dina(n3813), .dinb(n3804), .dout(n3814));
  jand g3173(.dina(n2628), .dinb(\in0[91] ), .dout(n3815));
  jand g3174(.dina(n2783), .dinb(\in1[91] ), .dout(n3816));
  jor  g3175(.dina(n3816), .dinb(n3815), .dout(n3817));
  jnot g3176(.din(n3817), .dout(n3818));
  jand g3177(.dina(n1556), .dinb(\in2[91] ), .dout(n3819));
  jand g3178(.dina(n1711), .dinb(\in3[91] ), .dout(n3820));
  jor  g3179(.dina(n3820), .dinb(n3819), .dout(n3821));
  jand g3180(.dina(n3821), .dinb(n3818), .dout(n3822));
  jand g3181(.dina(n1556), .dinb(\in2[90] ), .dout(n3823));
  jand g3182(.dina(n1711), .dinb(\in3[90] ), .dout(n3824));
  jor  g3183(.dina(n3824), .dinb(n3823), .dout(n3825));
  jand g3184(.dina(n2628), .dinb(\in0[90] ), .dout(n3826));
  jand g3185(.dina(n2783), .dinb(\in1[90] ), .dout(n3827));
  jor  g3186(.dina(n3827), .dinb(n3826), .dout(n3828));
  jnot g3187(.din(n3828), .dout(n3829));
  jand g3188(.dina(n3829), .dinb(n3825), .dout(n3830));
  jor  g3189(.dina(n3830), .dinb(n3822), .dout(n3831));
  jand g3190(.dina(n2628), .dinb(\in0[89] ), .dout(n3832));
  jand g3191(.dina(n2783), .dinb(\in1[89] ), .dout(n3833));
  jor  g3192(.dina(n3833), .dinb(n3832), .dout(n3834));
  jnot g3193(.din(n3834), .dout(n3835));
  jand g3194(.dina(n1556), .dinb(\in2[89] ), .dout(n3836));
  jand g3195(.dina(n1711), .dinb(\in3[89] ), .dout(n3837));
  jor  g3196(.dina(n3837), .dinb(n3836), .dout(n3838));
  jand g3197(.dina(n3838), .dinb(n3835), .dout(n3839));
  jand g3198(.dina(n1556), .dinb(\in2[88] ), .dout(n3840));
  jand g3199(.dina(n1711), .dinb(\in3[88] ), .dout(n3841));
  jor  g3200(.dina(n3841), .dinb(n3840), .dout(n3842));
  jand g3201(.dina(n2628), .dinb(\in0[88] ), .dout(n3843));
  jand g3202(.dina(n2783), .dinb(\in1[88] ), .dout(n3844));
  jor  g3203(.dina(n3844), .dinb(n3843), .dout(n3845));
  jnot g3204(.din(n3845), .dout(n3846));
  jand g3205(.dina(n3846), .dinb(n3842), .dout(n3847));
  jor  g3206(.dina(n3847), .dinb(n3839), .dout(n3848));
  jor  g3207(.dina(n3848), .dinb(n3831), .dout(n3849));
  jor  g3208(.dina(n3849), .dinb(n3814), .dout(n3850));
  jor  g3209(.dina(n3821), .dinb(n3818), .dout(n3851));
  jor  g3210(.dina(n3846), .dinb(n3842), .dout(n3852));
  jor  g3211(.dina(n3852), .dinb(n3839), .dout(n3853));
  jor  g3212(.dina(n3838), .dinb(n3835), .dout(n3854));
  jor  g3213(.dina(n3829), .dinb(n3825), .dout(n3855));
  jand g3214(.dina(n3855), .dinb(n3854), .dout(n3856));
  jand g3215(.dina(n3856), .dinb(n3853), .dout(n3857));
  jor  g3216(.dina(n3857), .dinb(n3831), .dout(n3858));
  jand g3217(.dina(n3858), .dinb(n3851), .dout(n3859));
  jand g3218(.dina(n3859), .dinb(n3850), .dout(n3860));
  jand g3219(.dina(n2628), .dinb(\in0[92] ), .dout(n3861));
  jand g3220(.dina(n2783), .dinb(\in1[92] ), .dout(n3862));
  jor  g3221(.dina(n3862), .dinb(n3861), .dout(n3863));
  jnot g3222(.din(n3863), .dout(n3864));
  jand g3223(.dina(n1556), .dinb(\in2[92] ), .dout(n3865));
  jand g3224(.dina(n1711), .dinb(\in3[92] ), .dout(n3866));
  jor  g3225(.dina(n3866), .dinb(n3865), .dout(n3867));
  jand g3226(.dina(n3867), .dinb(n3864), .dout(n3868));
  jand g3227(.dina(n2628), .dinb(\in0[93] ), .dout(n3869));
  jand g3228(.dina(n2783), .dinb(\in1[93] ), .dout(n3870));
  jor  g3229(.dina(n3870), .dinb(n3869), .dout(n3871));
  jnot g3230(.din(n3871), .dout(n3872));
  jand g3231(.dina(n1556), .dinb(\in2[93] ), .dout(n3873));
  jand g3232(.dina(n1711), .dinb(\in3[93] ), .dout(n3874));
  jor  g3233(.dina(n3874), .dinb(n3873), .dout(n3875));
  jand g3234(.dina(n3875), .dinb(n3872), .dout(n3876));
  jand g3235(.dina(n2628), .dinb(\in0[95] ), .dout(n3877));
  jand g3236(.dina(n2783), .dinb(\in1[95] ), .dout(n3878));
  jor  g3237(.dina(n3878), .dinb(n3877), .dout(n3879));
  jnot g3238(.din(n3879), .dout(n3880));
  jand g3239(.dina(n1556), .dinb(\in2[95] ), .dout(n3881));
  jand g3240(.dina(n1711), .dinb(\in3[95] ), .dout(n3882));
  jor  g3241(.dina(n3882), .dinb(n3881), .dout(n3883));
  jand g3242(.dina(n3883), .dinb(n3880), .dout(n3884));
  jand g3243(.dina(n1556), .dinb(\in2[94] ), .dout(n3885));
  jand g3244(.dina(n1711), .dinb(\in3[94] ), .dout(n3886));
  jor  g3245(.dina(n3886), .dinb(n3885), .dout(n3887));
  jand g3246(.dina(n2628), .dinb(\in0[94] ), .dout(n3888));
  jand g3247(.dina(n2783), .dinb(\in1[94] ), .dout(n3889));
  jor  g3248(.dina(n3889), .dinb(n3888), .dout(n3890));
  jnot g3249(.din(n3890), .dout(n3891));
  jand g3250(.dina(n3891), .dinb(n3887), .dout(n3892));
  jor  g3251(.dina(n3892), .dinb(n3884), .dout(n3893));
  jor  g3252(.dina(n3893), .dinb(n3876), .dout(n3894));
  jor  g3253(.dina(n3894), .dinb(n3868), .dout(n3895));
  jor  g3254(.dina(n3895), .dinb(n3860), .dout(n3896));
  jor  g3255(.dina(n3875), .dinb(n3872), .dout(n3897));
  jor  g3256(.dina(n3867), .dinb(n3864), .dout(n3898));
  jand g3257(.dina(n3898), .dinb(n3897), .dout(n3899));
  jor  g3258(.dina(n3899), .dinb(n3894), .dout(n3900));
  jor  g3259(.dina(n3883), .dinb(n3880), .dout(n3901));
  jor  g3260(.dina(n3891), .dinb(n3887), .dout(n3902));
  jor  g3261(.dina(n3902), .dinb(n3884), .dout(n3903));
  jand g3262(.dina(n3903), .dinb(n3901), .dout(n3904));
  jand g3263(.dina(n3904), .dinb(n3900), .dout(n3905));
  jand g3264(.dina(n3905), .dinb(n3896), .dout(n3906));
  jand g3265(.dina(n2628), .dinb(\in0[99] ), .dout(n3907));
  jand g3266(.dina(n2783), .dinb(\in1[99] ), .dout(n3908));
  jor  g3267(.dina(n3908), .dinb(n3907), .dout(n3909));
  jnot g3268(.din(n3909), .dout(n3910));
  jand g3269(.dina(n1556), .dinb(\in2[99] ), .dout(n3911));
  jand g3270(.dina(n1711), .dinb(\in3[99] ), .dout(n3912));
  jor  g3271(.dina(n3912), .dinb(n3911), .dout(n3913));
  jand g3272(.dina(n3913), .dinb(n3910), .dout(n3914));
  jand g3273(.dina(n1556), .dinb(\in2[98] ), .dout(n3915));
  jand g3274(.dina(n1711), .dinb(\in3[98] ), .dout(n3916));
  jor  g3275(.dina(n3916), .dinb(n3915), .dout(n3917));
  jand g3276(.dina(n2628), .dinb(\in0[98] ), .dout(n3918));
  jand g3277(.dina(n2783), .dinb(\in1[98] ), .dout(n3919));
  jor  g3278(.dina(n3919), .dinb(n3918), .dout(n3920));
  jnot g3279(.din(n3920), .dout(n3921));
  jand g3280(.dina(n3921), .dinb(n3917), .dout(n3922));
  jor  g3281(.dina(n3922), .dinb(n3914), .dout(n3923));
  jand g3282(.dina(n2628), .dinb(\in0[97] ), .dout(n3924));
  jand g3283(.dina(n2783), .dinb(\in1[97] ), .dout(n3925));
  jor  g3284(.dina(n3925), .dinb(n3924), .dout(n3926));
  jnot g3285(.din(n3926), .dout(n3927));
  jand g3286(.dina(n1556), .dinb(\in2[97] ), .dout(n3928));
  jand g3287(.dina(n1711), .dinb(\in3[97] ), .dout(n3929));
  jor  g3288(.dina(n3929), .dinb(n3928), .dout(n3930));
  jand g3289(.dina(n3930), .dinb(n3927), .dout(n3931));
  jand g3290(.dina(n1556), .dinb(\in2[96] ), .dout(n3932));
  jand g3291(.dina(n1711), .dinb(\in3[96] ), .dout(n3933));
  jor  g3292(.dina(n3933), .dinb(n3932), .dout(n3934));
  jand g3293(.dina(n2628), .dinb(\in0[96] ), .dout(n3935));
  jand g3294(.dina(n2783), .dinb(\in1[96] ), .dout(n3936));
  jor  g3295(.dina(n3936), .dinb(n3935), .dout(n3937));
  jnot g3296(.din(n3937), .dout(n3938));
  jand g3297(.dina(n3938), .dinb(n3934), .dout(n3939));
  jor  g3298(.dina(n3939), .dinb(n3931), .dout(n3940));
  jor  g3299(.dina(n3940), .dinb(n3923), .dout(n3941));
  jor  g3300(.dina(n3941), .dinb(n3906), .dout(n3942));
  jor  g3301(.dina(n3913), .dinb(n3910), .dout(n3943));
  jor  g3302(.dina(n3938), .dinb(n3934), .dout(n3944));
  jor  g3303(.dina(n3944), .dinb(n3931), .dout(n3945));
  jor  g3304(.dina(n3930), .dinb(n3927), .dout(n3946));
  jor  g3305(.dina(n3921), .dinb(n3917), .dout(n3947));
  jand g3306(.dina(n3947), .dinb(n3946), .dout(n3948));
  jand g3307(.dina(n3948), .dinb(n3945), .dout(n3949));
  jor  g3308(.dina(n3949), .dinb(n3923), .dout(n3950));
  jand g3309(.dina(n3950), .dinb(n3943), .dout(n3951));
  jand g3310(.dina(n3951), .dinb(n3942), .dout(n3952));
  jand g3311(.dina(n2628), .dinb(\in0[100] ), .dout(n3953));
  jand g3312(.dina(n2783), .dinb(\in1[100] ), .dout(n3954));
  jor  g3313(.dina(n3954), .dinb(n3953), .dout(n3955));
  jnot g3314(.din(n3955), .dout(n3956));
  jand g3315(.dina(n1556), .dinb(\in2[100] ), .dout(n3957));
  jand g3316(.dina(n1711), .dinb(\in3[100] ), .dout(n3958));
  jor  g3317(.dina(n3958), .dinb(n3957), .dout(n3959));
  jand g3318(.dina(n3959), .dinb(n3956), .dout(n3960));
  jand g3319(.dina(n2628), .dinb(\in0[101] ), .dout(n3961));
  jand g3320(.dina(n2783), .dinb(\in1[101] ), .dout(n3962));
  jor  g3321(.dina(n3962), .dinb(n3961), .dout(n3963));
  jnot g3322(.din(n3963), .dout(n3964));
  jand g3323(.dina(n1556), .dinb(\in2[101] ), .dout(n3965));
  jand g3324(.dina(n1711), .dinb(\in3[101] ), .dout(n3966));
  jor  g3325(.dina(n3966), .dinb(n3965), .dout(n3967));
  jand g3326(.dina(n3967), .dinb(n3964), .dout(n3968));
  jand g3327(.dina(n2628), .dinb(\in0[103] ), .dout(n3969));
  jand g3328(.dina(n2783), .dinb(\in1[103] ), .dout(n3970));
  jor  g3329(.dina(n3970), .dinb(n3969), .dout(n3971));
  jnot g3330(.din(n3971), .dout(n3972));
  jand g3331(.dina(n1556), .dinb(\in2[103] ), .dout(n3973));
  jand g3332(.dina(n1711), .dinb(\in3[103] ), .dout(n3974));
  jor  g3333(.dina(n3974), .dinb(n3973), .dout(n3975));
  jand g3334(.dina(n3975), .dinb(n3972), .dout(n3976));
  jand g3335(.dina(n1556), .dinb(\in2[102] ), .dout(n3977));
  jand g3336(.dina(n1711), .dinb(\in3[102] ), .dout(n3978));
  jor  g3337(.dina(n3978), .dinb(n3977), .dout(n3979));
  jand g3338(.dina(n2628), .dinb(\in0[102] ), .dout(n3980));
  jand g3339(.dina(n2783), .dinb(\in1[102] ), .dout(n3981));
  jor  g3340(.dina(n3981), .dinb(n3980), .dout(n3982));
  jnot g3341(.din(n3982), .dout(n3983));
  jand g3342(.dina(n3983), .dinb(n3979), .dout(n3984));
  jor  g3343(.dina(n3984), .dinb(n3976), .dout(n3985));
  jor  g3344(.dina(n3985), .dinb(n3968), .dout(n3986));
  jor  g3345(.dina(n3986), .dinb(n3960), .dout(n3987));
  jor  g3346(.dina(n3987), .dinb(n3952), .dout(n3988));
  jor  g3347(.dina(n3967), .dinb(n3964), .dout(n3989));
  jor  g3348(.dina(n3959), .dinb(n3956), .dout(n3990));
  jand g3349(.dina(n3990), .dinb(n3989), .dout(n3991));
  jor  g3350(.dina(n3991), .dinb(n3986), .dout(n3992));
  jor  g3351(.dina(n3975), .dinb(n3972), .dout(n3993));
  jor  g3352(.dina(n3983), .dinb(n3979), .dout(n3994));
  jor  g3353(.dina(n3994), .dinb(n3976), .dout(n3995));
  jand g3354(.dina(n3995), .dinb(n3993), .dout(n3996));
  jand g3355(.dina(n3996), .dinb(n3992), .dout(n3997));
  jand g3356(.dina(n3997), .dinb(n3988), .dout(n3998));
  jand g3357(.dina(n2628), .dinb(\in0[107] ), .dout(n3999));
  jand g3358(.dina(n2783), .dinb(\in1[107] ), .dout(n4000));
  jor  g3359(.dina(n4000), .dinb(n3999), .dout(n4001));
  jnot g3360(.din(n4001), .dout(n4002));
  jand g3361(.dina(n1556), .dinb(\in2[107] ), .dout(n4003));
  jand g3362(.dina(n1711), .dinb(\in3[107] ), .dout(n4004));
  jor  g3363(.dina(n4004), .dinb(n4003), .dout(n4005));
  jand g3364(.dina(n4005), .dinb(n4002), .dout(n4006));
  jand g3365(.dina(n1556), .dinb(\in2[106] ), .dout(n4007));
  jand g3366(.dina(n1711), .dinb(\in3[106] ), .dout(n4008));
  jor  g3367(.dina(n4008), .dinb(n4007), .dout(n4009));
  jand g3368(.dina(n2628), .dinb(\in0[106] ), .dout(n4010));
  jand g3369(.dina(n2783), .dinb(\in1[106] ), .dout(n4011));
  jor  g3370(.dina(n4011), .dinb(n4010), .dout(n4012));
  jnot g3371(.din(n4012), .dout(n4013));
  jand g3372(.dina(n4013), .dinb(n4009), .dout(n4014));
  jor  g3373(.dina(n4014), .dinb(n4006), .dout(n4015));
  jand g3374(.dina(n2628), .dinb(\in0[105] ), .dout(n4016));
  jand g3375(.dina(n2783), .dinb(\in1[105] ), .dout(n4017));
  jor  g3376(.dina(n4017), .dinb(n4016), .dout(n4018));
  jnot g3377(.din(n4018), .dout(n4019));
  jand g3378(.dina(n1556), .dinb(\in2[105] ), .dout(n4020));
  jand g3379(.dina(n1711), .dinb(\in3[105] ), .dout(n4021));
  jor  g3380(.dina(n4021), .dinb(n4020), .dout(n4022));
  jand g3381(.dina(n4022), .dinb(n4019), .dout(n4023));
  jand g3382(.dina(n1556), .dinb(\in2[104] ), .dout(n4024));
  jand g3383(.dina(n1711), .dinb(\in3[104] ), .dout(n4025));
  jor  g3384(.dina(n4025), .dinb(n4024), .dout(n4026));
  jand g3385(.dina(n2628), .dinb(\in0[104] ), .dout(n4027));
  jand g3386(.dina(n2783), .dinb(\in1[104] ), .dout(n4028));
  jor  g3387(.dina(n4028), .dinb(n4027), .dout(n4029));
  jnot g3388(.din(n4029), .dout(n4030));
  jand g3389(.dina(n4030), .dinb(n4026), .dout(n4031));
  jor  g3390(.dina(n4031), .dinb(n4023), .dout(n4032));
  jor  g3391(.dina(n4032), .dinb(n4015), .dout(n4033));
  jor  g3392(.dina(n4033), .dinb(n3998), .dout(n4034));
  jor  g3393(.dina(n4005), .dinb(n4002), .dout(n4035));
  jor  g3394(.dina(n4030), .dinb(n4026), .dout(n4036));
  jor  g3395(.dina(n4036), .dinb(n4023), .dout(n4037));
  jor  g3396(.dina(n4022), .dinb(n4019), .dout(n4038));
  jor  g3397(.dina(n4013), .dinb(n4009), .dout(n4039));
  jand g3398(.dina(n4039), .dinb(n4038), .dout(n4040));
  jand g3399(.dina(n4040), .dinb(n4037), .dout(n4041));
  jor  g3400(.dina(n4041), .dinb(n4015), .dout(n4042));
  jand g3401(.dina(n4042), .dinb(n4035), .dout(n4043));
  jand g3402(.dina(n4043), .dinb(n4034), .dout(n4044));
  jand g3403(.dina(n2628), .dinb(\in0[108] ), .dout(n4045));
  jand g3404(.dina(n2783), .dinb(\in1[108] ), .dout(n4046));
  jor  g3405(.dina(n4046), .dinb(n4045), .dout(n4047));
  jnot g3406(.din(n4047), .dout(n4048));
  jand g3407(.dina(n1556), .dinb(\in2[108] ), .dout(n4049));
  jand g3408(.dina(n1711), .dinb(\in3[108] ), .dout(n4050));
  jor  g3409(.dina(n4050), .dinb(n4049), .dout(n4051));
  jand g3410(.dina(n4051), .dinb(n4048), .dout(n4052));
  jand g3411(.dina(n2628), .dinb(\in0[109] ), .dout(n4053));
  jand g3412(.dina(n2783), .dinb(\in1[109] ), .dout(n4054));
  jor  g3413(.dina(n4054), .dinb(n4053), .dout(n4055));
  jnot g3414(.din(n4055), .dout(n4056));
  jand g3415(.dina(n1556), .dinb(\in2[109] ), .dout(n4057));
  jand g3416(.dina(n1711), .dinb(\in3[109] ), .dout(n4058));
  jor  g3417(.dina(n4058), .dinb(n4057), .dout(n4059));
  jand g3418(.dina(n4059), .dinb(n4056), .dout(n4060));
  jand g3419(.dina(n2628), .dinb(\in0[111] ), .dout(n4061));
  jand g3420(.dina(n2783), .dinb(\in1[111] ), .dout(n4062));
  jor  g3421(.dina(n4062), .dinb(n4061), .dout(n4063));
  jnot g3422(.din(n4063), .dout(n4064));
  jand g3423(.dina(n1556), .dinb(\in2[111] ), .dout(n4065));
  jand g3424(.dina(n1711), .dinb(\in3[111] ), .dout(n4066));
  jor  g3425(.dina(n4066), .dinb(n4065), .dout(n4067));
  jand g3426(.dina(n4067), .dinb(n4064), .dout(n4068));
  jand g3427(.dina(n1556), .dinb(\in2[110] ), .dout(n4069));
  jand g3428(.dina(n1711), .dinb(\in3[110] ), .dout(n4070));
  jor  g3429(.dina(n4070), .dinb(n4069), .dout(n4071));
  jand g3430(.dina(n2628), .dinb(\in0[110] ), .dout(n4072));
  jand g3431(.dina(n2783), .dinb(\in1[110] ), .dout(n4073));
  jor  g3432(.dina(n4073), .dinb(n4072), .dout(n4074));
  jnot g3433(.din(n4074), .dout(n4075));
  jand g3434(.dina(n4075), .dinb(n4071), .dout(n4076));
  jor  g3435(.dina(n4076), .dinb(n4068), .dout(n4077));
  jor  g3436(.dina(n4077), .dinb(n4060), .dout(n4078));
  jor  g3437(.dina(n4078), .dinb(n4052), .dout(n4079));
  jor  g3438(.dina(n4079), .dinb(n4044), .dout(n4080));
  jor  g3439(.dina(n4059), .dinb(n4056), .dout(n4081));
  jor  g3440(.dina(n4051), .dinb(n4048), .dout(n4082));
  jand g3441(.dina(n4082), .dinb(n4081), .dout(n4083));
  jor  g3442(.dina(n4083), .dinb(n4078), .dout(n4084));
  jor  g3443(.dina(n4067), .dinb(n4064), .dout(n4085));
  jor  g3444(.dina(n4075), .dinb(n4071), .dout(n4086));
  jor  g3445(.dina(n4086), .dinb(n4068), .dout(n4087));
  jand g3446(.dina(n4087), .dinb(n4085), .dout(n4088));
  jand g3447(.dina(n4088), .dinb(n4084), .dout(n4089));
  jand g3448(.dina(n4089), .dinb(n4080), .dout(n4090));
  jand g3449(.dina(n2628), .dinb(\in0[115] ), .dout(n4091));
  jand g3450(.dina(n2783), .dinb(\in1[115] ), .dout(n4092));
  jor  g3451(.dina(n4092), .dinb(n4091), .dout(n4093));
  jnot g3452(.din(n4093), .dout(n4094));
  jand g3453(.dina(n1556), .dinb(\in2[115] ), .dout(n4095));
  jand g3454(.dina(n1711), .dinb(\in3[115] ), .dout(n4096));
  jor  g3455(.dina(n4096), .dinb(n4095), .dout(n4097));
  jand g3456(.dina(n4097), .dinb(n4094), .dout(n4098));
  jand g3457(.dina(n1556), .dinb(\in2[114] ), .dout(n4099));
  jand g3458(.dina(n1711), .dinb(\in3[114] ), .dout(n4100));
  jor  g3459(.dina(n4100), .dinb(n4099), .dout(n4101));
  jand g3460(.dina(n2628), .dinb(\in0[114] ), .dout(n4102));
  jand g3461(.dina(n2783), .dinb(\in1[114] ), .dout(n4103));
  jor  g3462(.dina(n4103), .dinb(n4102), .dout(n4104));
  jnot g3463(.din(n4104), .dout(n4105));
  jand g3464(.dina(n4105), .dinb(n4101), .dout(n4106));
  jor  g3465(.dina(n4106), .dinb(n4098), .dout(n4107));
  jand g3466(.dina(n2628), .dinb(\in0[113] ), .dout(n4108));
  jand g3467(.dina(n2783), .dinb(\in1[113] ), .dout(n4109));
  jor  g3468(.dina(n4109), .dinb(n4108), .dout(n4110));
  jnot g3469(.din(n4110), .dout(n4111));
  jand g3470(.dina(n1556), .dinb(\in2[113] ), .dout(n4112));
  jand g3471(.dina(n1711), .dinb(\in3[113] ), .dout(n4113));
  jor  g3472(.dina(n4113), .dinb(n4112), .dout(n4114));
  jand g3473(.dina(n4114), .dinb(n4111), .dout(n4115));
  jand g3474(.dina(n1556), .dinb(\in2[112] ), .dout(n4116));
  jand g3475(.dina(n1711), .dinb(\in3[112] ), .dout(n4117));
  jor  g3476(.dina(n4117), .dinb(n4116), .dout(n4118));
  jand g3477(.dina(n2628), .dinb(\in0[112] ), .dout(n4119));
  jand g3478(.dina(n2783), .dinb(\in1[112] ), .dout(n4120));
  jor  g3479(.dina(n4120), .dinb(n4119), .dout(n4121));
  jnot g3480(.din(n4121), .dout(n4122));
  jand g3481(.dina(n4122), .dinb(n4118), .dout(n4123));
  jor  g3482(.dina(n4123), .dinb(n4115), .dout(n4124));
  jor  g3483(.dina(n4124), .dinb(n4107), .dout(n4125));
  jor  g3484(.dina(n4125), .dinb(n4090), .dout(n4126));
  jor  g3485(.dina(n4097), .dinb(n4094), .dout(n4127));
  jor  g3486(.dina(n4122), .dinb(n4118), .dout(n4128));
  jor  g3487(.dina(n4128), .dinb(n4115), .dout(n4129));
  jor  g3488(.dina(n4114), .dinb(n4111), .dout(n4130));
  jor  g3489(.dina(n4105), .dinb(n4101), .dout(n4131));
  jand g3490(.dina(n4131), .dinb(n4130), .dout(n4132));
  jand g3491(.dina(n4132), .dinb(n4129), .dout(n4133));
  jor  g3492(.dina(n4133), .dinb(n4107), .dout(n4134));
  jand g3493(.dina(n4134), .dinb(n4127), .dout(n4135));
  jand g3494(.dina(n4135), .dinb(n4126), .dout(n4136));
  jand g3495(.dina(n2628), .dinb(\in0[116] ), .dout(n4137));
  jand g3496(.dina(n2783), .dinb(\in1[116] ), .dout(n4138));
  jor  g3497(.dina(n4138), .dinb(n4137), .dout(n4139));
  jnot g3498(.din(n4139), .dout(n4140));
  jand g3499(.dina(n1556), .dinb(\in2[116] ), .dout(n4141));
  jand g3500(.dina(n1711), .dinb(\in3[116] ), .dout(n4142));
  jor  g3501(.dina(n4142), .dinb(n4141), .dout(n4143));
  jand g3502(.dina(n4143), .dinb(n4140), .dout(n4144));
  jand g3503(.dina(n2628), .dinb(\in0[117] ), .dout(n4145));
  jand g3504(.dina(n2783), .dinb(\in1[117] ), .dout(n4146));
  jor  g3505(.dina(n4146), .dinb(n4145), .dout(n4147));
  jnot g3506(.din(n4147), .dout(n4148));
  jand g3507(.dina(n1556), .dinb(\in2[117] ), .dout(n4149));
  jand g3508(.dina(n1711), .dinb(\in3[117] ), .dout(n4150));
  jor  g3509(.dina(n4150), .dinb(n4149), .dout(n4151));
  jand g3510(.dina(n4151), .dinb(n4148), .dout(n4152));
  jand g3511(.dina(n2628), .dinb(\in0[119] ), .dout(n4153));
  jand g3512(.dina(n2783), .dinb(\in1[119] ), .dout(n4154));
  jor  g3513(.dina(n4154), .dinb(n4153), .dout(n4155));
  jnot g3514(.din(n4155), .dout(n4156));
  jand g3515(.dina(n1556), .dinb(\in2[119] ), .dout(n4157));
  jand g3516(.dina(n1711), .dinb(\in3[119] ), .dout(n4158));
  jor  g3517(.dina(n4158), .dinb(n4157), .dout(n4159));
  jand g3518(.dina(n4159), .dinb(n4156), .dout(n4160));
  jand g3519(.dina(n1556), .dinb(\in2[118] ), .dout(n4161));
  jand g3520(.dina(n1711), .dinb(\in3[118] ), .dout(n4162));
  jor  g3521(.dina(n4162), .dinb(n4161), .dout(n4163));
  jand g3522(.dina(n2628), .dinb(\in0[118] ), .dout(n4164));
  jand g3523(.dina(n2783), .dinb(\in1[118] ), .dout(n4165));
  jor  g3524(.dina(n4165), .dinb(n4164), .dout(n4166));
  jnot g3525(.din(n4166), .dout(n4167));
  jand g3526(.dina(n4167), .dinb(n4163), .dout(n4168));
  jor  g3527(.dina(n4168), .dinb(n4160), .dout(n4169));
  jor  g3528(.dina(n4169), .dinb(n4152), .dout(n4170));
  jor  g3529(.dina(n4170), .dinb(n4144), .dout(n4171));
  jor  g3530(.dina(n4171), .dinb(n4136), .dout(n4172));
  jor  g3531(.dina(n4151), .dinb(n4148), .dout(n4173));
  jor  g3532(.dina(n4143), .dinb(n4140), .dout(n4174));
  jand g3533(.dina(n4174), .dinb(n4173), .dout(n4175));
  jor  g3534(.dina(n4175), .dinb(n4170), .dout(n4176));
  jor  g3535(.dina(n4159), .dinb(n4156), .dout(n4177));
  jor  g3536(.dina(n4167), .dinb(n4163), .dout(n4178));
  jor  g3537(.dina(n4178), .dinb(n4160), .dout(n4179));
  jand g3538(.dina(n4179), .dinb(n4177), .dout(n4180));
  jand g3539(.dina(n4180), .dinb(n4176), .dout(n4181));
  jand g3540(.dina(n4181), .dinb(n4172), .dout(n4182));
  jand g3541(.dina(n2628), .dinb(\in0[123] ), .dout(n4183));
  jand g3542(.dina(n2783), .dinb(\in1[123] ), .dout(n4184));
  jor  g3543(.dina(n4184), .dinb(n4183), .dout(n4185));
  jnot g3544(.din(n4185), .dout(n4186));
  jand g3545(.dina(n1556), .dinb(\in2[123] ), .dout(n4187));
  jand g3546(.dina(n1711), .dinb(\in3[123] ), .dout(n4188));
  jor  g3547(.dina(n4188), .dinb(n4187), .dout(n4189));
  jand g3548(.dina(n4189), .dinb(n4186), .dout(n4190));
  jand g3549(.dina(n1556), .dinb(\in2[122] ), .dout(n4191));
  jand g3550(.dina(n1711), .dinb(\in3[122] ), .dout(n4192));
  jor  g3551(.dina(n4192), .dinb(n4191), .dout(n4193));
  jand g3552(.dina(n2628), .dinb(\in0[122] ), .dout(n4194));
  jand g3553(.dina(n2783), .dinb(\in1[122] ), .dout(n4195));
  jor  g3554(.dina(n4195), .dinb(n4194), .dout(n4196));
  jnot g3555(.din(n4196), .dout(n4197));
  jand g3556(.dina(n4197), .dinb(n4193), .dout(n4198));
  jor  g3557(.dina(n4198), .dinb(n4190), .dout(n4199));
  jand g3558(.dina(n2628), .dinb(\in0[121] ), .dout(n4200));
  jand g3559(.dina(n2783), .dinb(\in1[121] ), .dout(n4201));
  jor  g3560(.dina(n4201), .dinb(n4200), .dout(n4202));
  jnot g3561(.din(n4202), .dout(n4203));
  jand g3562(.dina(n1556), .dinb(\in2[121] ), .dout(n4204));
  jand g3563(.dina(n1711), .dinb(\in3[121] ), .dout(n4205));
  jor  g3564(.dina(n4205), .dinb(n4204), .dout(n4206));
  jand g3565(.dina(n4206), .dinb(n4203), .dout(n4207));
  jand g3566(.dina(n1556), .dinb(\in2[120] ), .dout(n4208));
  jand g3567(.dina(n1711), .dinb(\in3[120] ), .dout(n4209));
  jor  g3568(.dina(n4209), .dinb(n4208), .dout(n4210));
  jand g3569(.dina(n2628), .dinb(\in0[120] ), .dout(n4211));
  jand g3570(.dina(n2783), .dinb(\in1[120] ), .dout(n4212));
  jor  g3571(.dina(n4212), .dinb(n4211), .dout(n4213));
  jnot g3572(.din(n4213), .dout(n4214));
  jand g3573(.dina(n4214), .dinb(n4210), .dout(n4215));
  jor  g3574(.dina(n4215), .dinb(n4207), .dout(n4216));
  jor  g3575(.dina(n4216), .dinb(n4199), .dout(n4217));
  jor  g3576(.dina(n4217), .dinb(n4182), .dout(n4218));
  jor  g3577(.dina(n4189), .dinb(n4186), .dout(n4219));
  jor  g3578(.dina(n4214), .dinb(n4210), .dout(n4220));
  jor  g3579(.dina(n4220), .dinb(n4207), .dout(n4221));
  jor  g3580(.dina(n4206), .dinb(n4203), .dout(n4222));
  jor  g3581(.dina(n4197), .dinb(n4193), .dout(n4223));
  jand g3582(.dina(n4223), .dinb(n4222), .dout(n4224));
  jand g3583(.dina(n4224), .dinb(n4221), .dout(n4225));
  jor  g3584(.dina(n4225), .dinb(n4199), .dout(n4226));
  jand g3585(.dina(n4226), .dinb(n4219), .dout(n4227));
  jand g3586(.dina(n4227), .dinb(n4218), .dout(n4228));
  jand g3587(.dina(n2628), .dinb(\in0[126] ), .dout(n4229));
  jand g3588(.dina(n2783), .dinb(\in1[126] ), .dout(n4230));
  jor  g3589(.dina(n4230), .dinb(n4229), .dout(n4231));
  jnot g3590(.din(n4231), .dout(n4232));
  jand g3591(.dina(n1556), .dinb(\in2[126] ), .dout(n4233));
  jand g3592(.dina(n1711), .dinb(\in3[126] ), .dout(n4234));
  jor  g3593(.dina(n4234), .dinb(n4233), .dout(n4235));
  jand g3594(.dina(n4235), .dinb(n4232), .dout(n4236));
  jand g3595(.dina(n2628), .dinb(\in0[125] ), .dout(n4237));
  jand g3596(.dina(n2783), .dinb(\in1[125] ), .dout(n4238));
  jor  g3597(.dina(n4238), .dinb(n4237), .dout(n4239));
  jnot g3598(.din(n4239), .dout(n4240));
  jand g3599(.dina(n1556), .dinb(\in2[125] ), .dout(n4241));
  jand g3600(.dina(n1711), .dinb(\in3[125] ), .dout(n4242));
  jor  g3601(.dina(n4242), .dinb(n4241), .dout(n4243));
  jand g3602(.dina(n4243), .dinb(n4240), .dout(n4244));
  jor  g3603(.dina(n4244), .dinb(n4236), .dout(n4245));
  jand g3604(.dina(\in3[127] ), .dinb(\in2[127] ), .dout(n4246));
  jnot g3605(.din(n4246), .dout(n4247));
  jand g3606(.dina(\in1[127] ), .dinb(\in0[127] ), .dout(n4248));
  jand g3607(.dina(n4248), .dinb(n4247), .dout(n4249));
  jand g3608(.dina(n2628), .dinb(\in0[124] ), .dout(n4250));
  jand g3609(.dina(n2783), .dinb(\in1[124] ), .dout(n4251));
  jor  g3610(.dina(n4251), .dinb(n4250), .dout(n4252));
  jnot g3611(.din(n4252), .dout(n4253));
  jand g3612(.dina(n1556), .dinb(\in2[124] ), .dout(n4254));
  jand g3613(.dina(n1711), .dinb(\in3[124] ), .dout(n4255));
  jor  g3614(.dina(n4255), .dinb(n4254), .dout(n4256));
  jand g3615(.dina(n4256), .dinb(n4253), .dout(n4257));
  jor  g3616(.dina(n4257), .dinb(n4249), .dout(n4258));
  jor  g3617(.dina(n4258), .dinb(n4245), .dout(n4259));
  jor  g3618(.dina(n4259), .dinb(n4228), .dout(n4260));
  jor  g3619(.dina(n4256), .dinb(n4253), .dout(n4261));
  jor  g3620(.dina(n4243), .dinb(n4240), .dout(n4262));
  jand g3621(.dina(n4262), .dinb(n4261), .dout(n4263));
  jor  g3622(.dina(n4263), .dinb(n4245), .dout(n4264));
  jor  g3623(.dina(n4248), .dinb(n4247), .dout(n4265));
  jor  g3624(.dina(n4235), .dinb(n4232), .dout(n4266));
  jand g3625(.dina(n4266), .dinb(n4265), .dout(n4267));
  jand g3626(.dina(n4267), .dinb(n4264), .dout(n4268));
  jor  g3627(.dina(n4268), .dinb(n4249), .dout(n4269));
  jand g3628(.dina(n4269), .dinb(n4260), .dout(\address[1] ));
  jand g3629(.dina(\address[1] ), .dinb(n1713), .dout(n4271));
  jand g3630(.dina(n2628), .dinb(\in0[0] ), .dout(n4272));
  jand g3631(.dina(n2783), .dinb(\in1[0] ), .dout(n4273));
  jor  g3632(.dina(n4273), .dinb(n4272), .dout(n4274));
  jnot g3633(.din(n2790), .dout(n4275));
  jnot g3634(.din(n2862), .dout(n4276));
  jnot g3635(.din(n2896), .dout(n4277));
  jnot g3636(.din(n2908), .dout(n4278));
  jnot g3637(.din(n2909), .dout(n4279));
  jnot g3638(.din(n2917), .dout(n4280));
  jnot g3639(.din(n2925), .dout(n4281));
  jnot g3640(.din(n2983), .dout(n4282));
  jnot g3641(.din(n3010), .dout(n4283));
  jnot g3642(.din(n3011), .dout(n4284));
  jnot g3643(.din(n3018), .dout(n4285));
  jnot g3644(.din(n3021), .dout(n4286));
  jor  g3645(.dina(n1711), .dinb(n1589), .dout(n4287));
  jor  g3646(.dina(n1556), .dinb(n788), .dout(n4288));
  jand g3647(.dina(n4288), .dinb(n4287), .dout(n4289));
  jand g3648(.dina(n4274), .dinb(n4289), .dout(n4290));
  jand g3649(.dina(n2628), .dinb(\in0[1] ), .dout(n4291));
  jand g3650(.dina(n2783), .dinb(\in1[1] ), .dout(n4292));
  jor  g3651(.dina(n4292), .dinb(n4291), .dout(n4293));
  jor  g3652(.dina(n4293), .dinb(n4290), .dout(n4294));
  jand g3653(.dina(n4294), .dinb(n4286), .dout(n4295));
  jand g3654(.dina(n2628), .dinb(\in0[2] ), .dout(n4296));
  jand g3655(.dina(n2783), .dinb(\in1[2] ), .dout(n4297));
  jor  g3656(.dina(n4297), .dinb(n4296), .dout(n4298));
  jor  g3657(.dina(n1711), .dinb(n782), .dout(n4299));
  jor  g3658(.dina(n1556), .dinb(n780), .dout(n4300));
  jand g3659(.dina(n4300), .dinb(n4299), .dout(n4301));
  jand g3660(.dina(n4301), .dinb(n4298), .dout(n4302));
  jand g3661(.dina(n4293), .dinb(n4290), .dout(n4303));
  jor  g3662(.dina(n4303), .dinb(n4302), .dout(n4304));
  jor  g3663(.dina(n4304), .dinb(n4295), .dout(n4305));
  jand g3664(.dina(n4305), .dinb(n4285), .dout(n4306));
  jor  g3665(.dina(n4306), .dinb(n4284), .dout(n4307));
  jand g3666(.dina(n4307), .dinb(n4283), .dout(n4308));
  jnot g3667(.din(n3040), .dout(n4309));
  jand g3668(.dina(n4309), .dinb(n4308), .dout(n4310));
  jor  g3669(.dina(n4310), .dinb(n3001), .dout(n4311));
  jor  g3670(.dina(n4309), .dinb(n4308), .dout(n4312));
  jand g3671(.dina(n4312), .dinb(n4311), .dout(n4313));
  jnot g3672(.din(n3047), .dout(n4314));
  jand g3673(.dina(n4314), .dinb(n4313), .dout(n4315));
  jor  g3674(.dina(n4315), .dinb(n2997), .dout(n4316));
  jor  g3675(.dina(n4314), .dinb(n4313), .dout(n4317));
  jnot g3676(.din(n3058), .dout(n4318));
  jand g3677(.dina(n4318), .dinb(n4317), .dout(n4319));
  jand g3678(.dina(n4319), .dinb(n4316), .dout(n4320));
  jnot g3679(.din(n3061), .dout(n4321));
  jor  g3680(.dina(n4321), .dinb(n4320), .dout(n4322));
  jand g3681(.dina(n4322), .dinb(n2993), .dout(n4323));
  jor  g3682(.dina(n4323), .dinb(n2991), .dout(n4324));
  jor  g3683(.dina(n3067), .dinb(n4324), .dout(n4325));
  jand g3684(.dina(n4325), .dinb(n4282), .dout(n4326));
  jand g3685(.dina(n3067), .dinb(n4324), .dout(n4327));
  jor  g3686(.dina(n4327), .dinb(n4326), .dout(n4328));
  jand g3687(.dina(n4328), .dinb(n2979), .dout(n4329));
  jor  g3688(.dina(n4329), .dinb(n2977), .dout(n4330));
  jand g3689(.dina(n4330), .dinb(n2968), .dout(n4331));
  jor  g3690(.dina(n4331), .dinb(n2966), .dout(n4332));
  jand g3691(.dina(n4332), .dinb(n2957), .dout(n4333));
  jor  g3692(.dina(n4333), .dinb(n2955), .dout(n4334));
  jand g3693(.dina(n4334), .dinb(n2946), .dout(n4335));
  jor  g3694(.dina(n4335), .dinb(n2944), .dout(n4336));
  jand g3695(.dina(n4336), .dinb(n2935), .dout(n4337));
  jor  g3696(.dina(n4337), .dinb(n2933), .dout(n4338));
  jand g3697(.dina(n4338), .dinb(n4281), .dout(n4339));
  jnot g3698(.din(n3086), .dout(n4340));
  jor  g3699(.dina(n4340), .dinb(n4339), .dout(n4341));
  jand g3700(.dina(n4341), .dinb(n4280), .dout(n4342));
  jor  g3701(.dina(n4342), .dinb(n4279), .dout(n4343));
  jand g3702(.dina(n4343), .dinb(n4278), .dout(n4344));
  jor  g3703(.dina(n4344), .dinb(n2899), .dout(n4345));
  jand g3704(.dina(n4345), .dinb(n4277), .dout(n4346));
  jand g3705(.dina(n4344), .dinb(n2899), .dout(n4347));
  jor  g3706(.dina(n4347), .dinb(n3100), .dout(n4348));
  jor  g3707(.dina(n4348), .dinb(n4346), .dout(n4349));
  jand g3708(.dina(n3107), .dinb(n4349), .dout(n4350));
  jor  g3709(.dina(n4350), .dinb(n2892), .dout(n4351));
  jand g3710(.dina(n4351), .dinb(n2883), .dout(n4352));
  jor  g3711(.dina(n4352), .dinb(n2881), .dout(n4353));
  jand g3712(.dina(n4353), .dinb(n2872), .dout(n4354));
  jor  g3713(.dina(n4354), .dinb(n2870), .dout(n4355));
  jand g3714(.dina(n4355), .dinb(n4276), .dout(n4356));
  jnot g3715(.din(n3126), .dout(n4357));
  jor  g3716(.dina(n4357), .dinb(n4356), .dout(n4358));
  jand g3717(.dina(n3130), .dinb(n4358), .dout(n4359));
  jor  g3718(.dina(n4359), .dinb(n2853), .dout(n4360));
  jand g3719(.dina(n4360), .dinb(n2844), .dout(n4361));
  jor  g3720(.dina(n4361), .dinb(n2842), .dout(n4362));
  jand g3721(.dina(n4362), .dinb(n2833), .dout(n4363));
  jor  g3722(.dina(n4363), .dinb(n2831), .dout(n4364));
  jand g3723(.dina(n4364), .dinb(n2822), .dout(n4365));
  jor  g3724(.dina(n4365), .dinb(n2820), .dout(n4366));
  jand g3725(.dina(n4366), .dinb(n2811), .dout(n4367));
  jor  g3726(.dina(n4367), .dinb(n2809), .dout(n4368));
  jand g3727(.dina(n4368), .dinb(n2800), .dout(n4369));
  jor  g3728(.dina(n4369), .dinb(n2798), .dout(n4370));
  jand g3729(.dina(n4370), .dinb(n4275), .dout(n4371));
  jnot g3730(.din(n3155), .dout(n4372));
  jor  g3731(.dina(n4372), .dinb(n4371), .dout(n4373));
  jand g3732(.dina(n3233), .dinb(n4373), .dout(n4374));
  jnot g3733(.din(n3255), .dout(n4375));
  jor  g3734(.dina(n4375), .dinb(n4374), .dout(n4376));
  jnot g3735(.din(n3327), .dout(n4377));
  jand g3736(.dina(n4377), .dinb(n4376), .dout(n4378));
  jnot g3737(.din(n3348), .dout(n4379));
  jor  g3738(.dina(n4379), .dinb(n4378), .dout(n4380));
  jnot g3739(.din(n3423), .dout(n4381));
  jand g3740(.dina(n4381), .dinb(n4380), .dout(n4382));
  jnot g3741(.din(n3444), .dout(n4383));
  jor  g3742(.dina(n4383), .dinb(n4382), .dout(n4384));
  jnot g3743(.din(n3516), .dout(n4385));
  jand g3744(.dina(n4385), .dinb(n4384), .dout(n4386));
  jnot g3745(.din(n3537), .dout(n4387));
  jor  g3746(.dina(n4387), .dinb(n4386), .dout(n4388));
  jnot g3747(.din(n3573), .dout(n4389));
  jand g3748(.dina(n4389), .dinb(n4388), .dout(n4390));
  jnot g3749(.din(n3583), .dout(n4391));
  jor  g3750(.dina(n4391), .dinb(n4390), .dout(n4392));
  jnot g3751(.din(n3619), .dout(n4393));
  jand g3752(.dina(n4393), .dinb(n4392), .dout(n4394));
  jnot g3753(.din(n3629), .dout(n4395));
  jor  g3754(.dina(n4395), .dinb(n4394), .dout(n4396));
  jnot g3755(.din(n3665), .dout(n4397));
  jand g3756(.dina(n4397), .dinb(n4396), .dout(n4398));
  jnot g3757(.din(n3675), .dout(n4399));
  jor  g3758(.dina(n4399), .dinb(n4398), .dout(n4400));
  jnot g3759(.din(n3711), .dout(n4401));
  jand g3760(.dina(n4401), .dinb(n4400), .dout(n4402));
  jnot g3761(.din(n3721), .dout(n4403));
  jor  g3762(.dina(n4403), .dinb(n4402), .dout(n4404));
  jnot g3763(.din(n3757), .dout(n4405));
  jand g3764(.dina(n4405), .dinb(n4404), .dout(n4406));
  jnot g3765(.din(n3767), .dout(n4407));
  jor  g3766(.dina(n4407), .dinb(n4406), .dout(n4408));
  jnot g3767(.din(n3803), .dout(n4409));
  jand g3768(.dina(n4409), .dinb(n4408), .dout(n4410));
  jnot g3769(.din(n3813), .dout(n4411));
  jor  g3770(.dina(n4411), .dinb(n4410), .dout(n4412));
  jnot g3771(.din(n3849), .dout(n4413));
  jand g3772(.dina(n4413), .dinb(n4412), .dout(n4414));
  jnot g3773(.din(n3859), .dout(n4415));
  jor  g3774(.dina(n4415), .dinb(n4414), .dout(n4416));
  jnot g3775(.din(n3895), .dout(n4417));
  jand g3776(.dina(n4417), .dinb(n4416), .dout(n4418));
  jnot g3777(.din(n3905), .dout(n4419));
  jor  g3778(.dina(n4419), .dinb(n4418), .dout(n4420));
  jnot g3779(.din(n3941), .dout(n4421));
  jand g3780(.dina(n4421), .dinb(n4420), .dout(n4422));
  jnot g3781(.din(n3951), .dout(n4423));
  jor  g3782(.dina(n4423), .dinb(n4422), .dout(n4424));
  jnot g3783(.din(n3987), .dout(n4425));
  jand g3784(.dina(n4425), .dinb(n4424), .dout(n4426));
  jnot g3785(.din(n3997), .dout(n4427));
  jor  g3786(.dina(n4427), .dinb(n4426), .dout(n4428));
  jnot g3787(.din(n4033), .dout(n4429));
  jand g3788(.dina(n4429), .dinb(n4428), .dout(n4430));
  jnot g3789(.din(n4043), .dout(n4431));
  jor  g3790(.dina(n4431), .dinb(n4430), .dout(n4432));
  jnot g3791(.din(n4079), .dout(n4433));
  jand g3792(.dina(n4433), .dinb(n4432), .dout(n4434));
  jnot g3793(.din(n4089), .dout(n4435));
  jor  g3794(.dina(n4435), .dinb(n4434), .dout(n4436));
  jnot g3795(.din(n4125), .dout(n4437));
  jand g3796(.dina(n4437), .dinb(n4436), .dout(n4438));
  jnot g3797(.din(n4135), .dout(n4439));
  jor  g3798(.dina(n4439), .dinb(n4438), .dout(n4440));
  jnot g3799(.din(n4171), .dout(n4441));
  jand g3800(.dina(n4441), .dinb(n4440), .dout(n4442));
  jnot g3801(.din(n4181), .dout(n4443));
  jor  g3802(.dina(n4443), .dinb(n4442), .dout(n4444));
  jnot g3803(.din(n4217), .dout(n4445));
  jand g3804(.dina(n4445), .dinb(n4444), .dout(n4446));
  jnot g3805(.din(n4227), .dout(n4447));
  jor  g3806(.dina(n4447), .dinb(n4446), .dout(n4448));
  jnot g3807(.din(n4259), .dout(n4449));
  jand g3808(.dina(n4449), .dinb(n4448), .dout(n4450));
  jnot g3809(.din(n4269), .dout(n4451));
  jor  g3810(.dina(n4451), .dinb(n4450), .dout(n4452));
  jand g3811(.dina(n4452), .dinb(n4274), .dout(n4453));
  jor  g3812(.dina(n4453), .dinb(n4271), .dout(\result[0] ));
  jor  g3813(.dina(\address[1] ), .dinb(n4293), .dout(n4455));
  jor  g3814(.dina(n4452), .dinb(n3021), .dout(n4456));
  jand g3815(.dina(n4456), .dinb(n4455), .dout(\result[1] ));
  jor  g3816(.dina(\address[1] ), .dinb(n4298), .dout(n4458));
  jor  g3817(.dina(n4452), .dinb(n3017), .dout(n4459));
  jand g3818(.dina(n4459), .dinb(n4458), .dout(\result[2] ));
  jor  g3819(.dina(\address[1] ), .dinb(n3005), .dout(n4461));
  jor  g3820(.dina(n4452), .dinb(n3009), .dout(n4462));
  jand g3821(.dina(n4462), .dinb(n4461), .dout(\result[3] ));
  jand g3822(.dina(\address[1] ), .dinb(n3040), .dout(n4464));
  jand g3823(.dina(n4452), .dinb(n3001), .dout(n4465));
  jor  g3824(.dina(n4465), .dinb(n4464), .dout(\result[4] ));
  jand g3825(.dina(\address[1] ), .dinb(n3047), .dout(n4467));
  jand g3826(.dina(n4452), .dinb(n2997), .dout(n4468));
  jor  g3827(.dina(n4468), .dinb(n4467), .dout(\result[5] ));
  jand g3828(.dina(\address[1] ), .dinb(n3057), .dout(n4470));
  jand g3829(.dina(n4452), .dinb(n3053), .dout(n4471));
  jor  g3830(.dina(n4471), .dinb(n4470), .dout(\result[6] ));
  jor  g3831(.dina(\address[1] ), .dinb(n2986), .dout(n4473));
  jor  g3832(.dina(n4452), .dinb(n2989), .dout(n4474));
  jand g3833(.dina(n4474), .dinb(n4473), .dout(\result[7] ));
  jand g3834(.dina(\address[1] ), .dinb(n2983), .dout(n4476));
  jand g3835(.dina(n4452), .dinb(n3067), .dout(n4477));
  jor  g3836(.dina(n4477), .dinb(n4476), .dout(\result[8] ));
  jor  g3837(.dina(\address[1] ), .dinb(n2972), .dout(n4479));
  jor  g3838(.dina(n4452), .dinb(n2975), .dout(n4480));
  jand g3839(.dina(n4480), .dinb(n4479), .dout(\result[9] ));
  jor  g3840(.dina(\address[1] ), .dinb(n2961), .dout(n4482));
  jor  g3841(.dina(n4452), .dinb(n2964), .dout(n4483));
  jand g3842(.dina(n4483), .dinb(n4482), .dout(\result[10] ));
  jor  g3843(.dina(\address[1] ), .dinb(n2950), .dout(n4485));
  jor  g3844(.dina(n4452), .dinb(n2953), .dout(n4486));
  jand g3845(.dina(n4486), .dinb(n4485), .dout(\result[11] ));
  jor  g3846(.dina(\address[1] ), .dinb(n2939), .dout(n4488));
  jor  g3847(.dina(n4452), .dinb(n2942), .dout(n4489));
  jand g3848(.dina(n4489), .dinb(n4488), .dout(\result[12] ));
  jor  g3849(.dina(\address[1] ), .dinb(n2928), .dout(n4491));
  jor  g3850(.dina(n4452), .dinb(n2931), .dout(n4492));
  jand g3851(.dina(n4492), .dinb(n4491), .dout(\result[13] ));
  jor  g3852(.dina(\address[1] ), .dinb(n2920), .dout(n4494));
  jor  g3853(.dina(n4452), .dinb(n2924), .dout(n4495));
  jand g3854(.dina(n4495), .dinb(n4494), .dout(\result[14] ));
  jor  g3855(.dina(\address[1] ), .dinb(n2912), .dout(n4497));
  jor  g3856(.dina(n4452), .dinb(n2916), .dout(n4498));
  jand g3857(.dina(n4498), .dinb(n4497), .dout(\result[15] ));
  jor  g3858(.dina(\address[1] ), .dinb(n2903), .dout(n4500));
  jor  g3859(.dina(n4452), .dinb(n2907), .dout(n4501));
  jand g3860(.dina(n4501), .dinb(n4500), .dout(\result[16] ));
  jor  g3861(.dina(\address[1] ), .dinb(n2899), .dout(n4503));
  jor  g3862(.dina(n4452), .dinb(n2896), .dout(n4504));
  jand g3863(.dina(n4504), .dinb(n4503), .dout(\result[17] ));
  jor  g3864(.dina(\address[1] ), .dinb(n3095), .dout(n4506));
  jor  g3865(.dina(n4452), .dinb(n3098), .dout(n4507));
  jand g3866(.dina(n4507), .dinb(n4506), .dout(\result[18] ));
  jor  g3867(.dina(\address[1] ), .dinb(n2887), .dout(n4509));
  jor  g3868(.dina(n4452), .dinb(n2890), .dout(n4510));
  jand g3869(.dina(n4510), .dinb(n4509), .dout(\result[19] ));
  jor  g3870(.dina(\address[1] ), .dinb(n2876), .dout(n4512));
  jor  g3871(.dina(n4452), .dinb(n2879), .dout(n4513));
  jand g3872(.dina(n4513), .dinb(n4512), .dout(\result[20] ));
  jor  g3873(.dina(\address[1] ), .dinb(n2865), .dout(n4515));
  jor  g3874(.dina(n4452), .dinb(n2868), .dout(n4516));
  jand g3875(.dina(n4516), .dinb(n4515), .dout(\result[21] ));
  jor  g3876(.dina(\address[1] ), .dinb(n2857), .dout(n4518));
  jor  g3877(.dina(n4452), .dinb(n2861), .dout(n4519));
  jand g3878(.dina(n4519), .dinb(n4518), .dout(\result[22] ));
  jor  g3879(.dina(\address[1] ), .dinb(n3119), .dout(n4521));
  jor  g3880(.dina(n4452), .dinb(n3122), .dout(n4522));
  jand g3881(.dina(n4522), .dinb(n4521), .dout(\result[23] ));
  jor  g3882(.dina(\address[1] ), .dinb(n2848), .dout(n4524));
  jor  g3883(.dina(n4452), .dinb(n2851), .dout(n4525));
  jand g3884(.dina(n4525), .dinb(n4524), .dout(\result[24] ));
  jor  g3885(.dina(\address[1] ), .dinb(n2837), .dout(n4527));
  jor  g3886(.dina(n4452), .dinb(n2840), .dout(n4528));
  jand g3887(.dina(n4528), .dinb(n4527), .dout(\result[25] ));
  jor  g3888(.dina(\address[1] ), .dinb(n2826), .dout(n4530));
  jor  g3889(.dina(n4452), .dinb(n2829), .dout(n4531));
  jand g3890(.dina(n4531), .dinb(n4530), .dout(\result[26] ));
  jor  g3891(.dina(\address[1] ), .dinb(n2815), .dout(n4533));
  jor  g3892(.dina(n4452), .dinb(n2818), .dout(n4534));
  jand g3893(.dina(n4534), .dinb(n4533), .dout(\result[27] ));
  jor  g3894(.dina(\address[1] ), .dinb(n2804), .dout(n4536));
  jor  g3895(.dina(n4452), .dinb(n2807), .dout(n4537));
  jand g3896(.dina(n4537), .dinb(n4536), .dout(\result[28] ));
  jor  g3897(.dina(\address[1] ), .dinb(n2793), .dout(n4539));
  jor  g3898(.dina(n4452), .dinb(n2796), .dout(n4540));
  jand g3899(.dina(n4540), .dinb(n4539), .dout(\result[29] ));
  jor  g3900(.dina(\address[1] ), .dinb(n2785), .dout(n4542));
  jor  g3901(.dina(n4452), .dinb(n2789), .dout(n4543));
  jand g3902(.dina(n4543), .dinb(n4542), .dout(\result[30] ));
  jor  g3903(.dina(\address[1] ), .dinb(n3148), .dout(n4545));
  jor  g3904(.dina(n4452), .dinb(n3151), .dout(n4546));
  jand g3905(.dina(n4546), .dinb(n4545), .dout(\result[31] ));
  jor  g3906(.dina(\address[1] ), .dinb(n3216), .dout(n4548));
  jor  g3907(.dina(n4452), .dinb(n3213), .dout(n4549));
  jand g3908(.dina(n4549), .dinb(n4548), .dout(\result[32] ));
  jor  g3909(.dina(\address[1] ), .dinb(n3194), .dout(n4551));
  jor  g3910(.dina(n4452), .dinb(n3198), .dout(n4552));
  jand g3911(.dina(n4552), .dinb(n4551), .dout(\result[33] ));
  jor  g3912(.dina(\address[1] ), .dinb(n3205), .dout(n4554));
  jor  g3913(.dina(n4452), .dinb(n3202), .dout(n4555));
  jand g3914(.dina(n4555), .dinb(n4554), .dout(\result[34] ));
  jor  g3915(.dina(\address[1] ), .dinb(n3186), .dout(n4557));
  jor  g3916(.dina(n4452), .dinb(n3190), .dout(n4558));
  jand g3917(.dina(n4558), .dinb(n4557), .dout(\result[35] ));
  jor  g3918(.dina(\address[1] ), .dinb(n3222), .dout(n4560));
  jor  g3919(.dina(n4452), .dinb(n3226), .dout(n4561));
  jand g3920(.dina(n4561), .dinb(n4560), .dout(\result[36] ));
  jor  g3921(.dina(\address[1] ), .dinb(n3159), .dout(n4563));
  jor  g3922(.dina(n4452), .dinb(n3163), .dout(n4564));
  jand g3923(.dina(n4564), .dinb(n4563), .dout(\result[37] ));
  jor  g3924(.dina(\address[1] ), .dinb(n3178), .dout(n4566));
  jor  g3925(.dina(n4452), .dinb(n3175), .dout(n4567));
  jand g3926(.dina(n4567), .dinb(n4566), .dout(\result[38] ));
  jor  g3927(.dina(\address[1] ), .dinb(n3167), .dout(n4569));
  jor  g3928(.dina(n4452), .dinb(n3171), .dout(n4570));
  jand g3929(.dina(n4570), .dinb(n4569), .dout(\result[39] ));
  jor  g3930(.dina(\address[1] ), .dinb(n3310), .dout(n4572));
  jor  g3931(.dina(n4452), .dinb(n3314), .dout(n4573));
  jand g3932(.dina(n4573), .dinb(n4572), .dout(\result[40] ));
  jor  g3933(.dina(\address[1] ), .dinb(n3318), .dout(n4575));
  jor  g3934(.dina(n4452), .dinb(n3322), .dout(n4576));
  jand g3935(.dina(n4576), .dinb(n4575), .dout(\result[41] ));
  jor  g3936(.dina(\address[1] ), .dinb(n3293), .dout(n4578));
  jor  g3937(.dina(n4452), .dinb(n3297), .dout(n4579));
  jand g3938(.dina(n4579), .dinb(n4578), .dout(\result[42] ));
  jor  g3939(.dina(\address[1] ), .dinb(n3285), .dout(n4581));
  jor  g3940(.dina(n4452), .dinb(n3289), .dout(n4582));
  jand g3941(.dina(n4582), .dinb(n4581), .dout(\result[43] ));
  jor  g3942(.dina(\address[1] ), .dinb(n3302), .dout(n4584));
  jor  g3943(.dina(n4452), .dinb(n3306), .dout(n4585));
  jand g3944(.dina(n4585), .dinb(n4584), .dout(\result[44] ));
  jor  g3945(.dina(\address[1] ), .dinb(n3259), .dout(n4587));
  jor  g3946(.dina(n4452), .dinb(n3263), .dout(n4588));
  jand g3947(.dina(n4588), .dinb(n4587), .dout(\result[45] ));
  jor  g3948(.dina(\address[1] ), .dinb(n3278), .dout(n4590));
  jor  g3949(.dina(n4452), .dinb(n3275), .dout(n4591));
  jand g3950(.dina(n4591), .dinb(n4590), .dout(\result[46] ));
  jor  g3951(.dina(\address[1] ), .dinb(n3267), .dout(n4593));
  jor  g3952(.dina(n4452), .dinb(n3271), .dout(n4594));
  jand g3953(.dina(n4594), .dinb(n4593), .dout(\result[47] ));
  jor  g3954(.dina(\address[1] ), .dinb(n3418), .dout(n4596));
  jor  g3955(.dina(n4452), .dinb(n3415), .dout(n4597));
  jand g3956(.dina(n4597), .dinb(n4596), .dout(\result[48] ));
  jor  g3957(.dina(\address[1] ), .dinb(n3360), .dout(n4599));
  jor  g3958(.dina(n4452), .dinb(n3364), .dout(n4600));
  jand g3959(.dina(n4600), .dinb(n4599), .dout(\result[49] ));
  jor  g3960(.dina(\address[1] ), .dinb(n3371), .dout(n4602));
  jor  g3961(.dina(n4452), .dinb(n3368), .dout(n4603));
  jand g3962(.dina(n4603), .dinb(n4602), .dout(\result[50] ));
  jor  g3963(.dina(\address[1] ), .dinb(n3352), .dout(n4605));
  jor  g3964(.dina(n4452), .dinb(n3356), .dout(n4606));
  jand g3965(.dina(n4606), .dinb(n4605), .dout(\result[51] ));
  jor  g3966(.dina(\address[1] ), .dinb(n3387), .dout(n4608));
  jor  g3967(.dina(n4452), .dinb(n3391), .dout(n4609));
  jand g3968(.dina(n4609), .dinb(n4608), .dout(\result[52] ));
  jor  g3969(.dina(\address[1] ), .dinb(n3378), .dout(n4611));
  jor  g3970(.dina(n4452), .dinb(n3382), .dout(n4612));
  jand g3971(.dina(n4612), .dinb(n4611), .dout(\result[53] ));
  jor  g3972(.dina(\address[1] ), .dinb(n3409), .dout(n4614));
  jor  g3973(.dina(n4452), .dinb(n3406), .dout(n4615));
  jand g3974(.dina(n4615), .dinb(n4614), .dout(\result[54] ));
  jor  g3975(.dina(\address[1] ), .dinb(n3398), .dout(n4617));
  jor  g3976(.dina(n4452), .dinb(n3402), .dout(n4618));
  jand g3977(.dina(n4618), .dinb(n4617), .dout(\result[55] ));
  jor  g3978(.dina(\address[1] ), .dinb(n3499), .dout(n4620));
  jor  g3979(.dina(n4452), .dinb(n3503), .dout(n4621));
  jand g3980(.dina(n4621), .dinb(n4620), .dout(\result[56] ));
  jor  g3981(.dina(\address[1] ), .dinb(n3507), .dout(n4623));
  jor  g3982(.dina(n4452), .dinb(n3511), .dout(n4624));
  jand g3983(.dina(n4624), .dinb(n4623), .dout(\result[57] ));
  jor  g3984(.dina(\address[1] ), .dinb(n3482), .dout(n4626));
  jor  g3985(.dina(n4452), .dinb(n3486), .dout(n4627));
  jand g3986(.dina(n4627), .dinb(n4626), .dout(\result[58] ));
  jor  g3987(.dina(\address[1] ), .dinb(n3474), .dout(n4629));
  jor  g3988(.dina(n4452), .dinb(n3478), .dout(n4630));
  jand g3989(.dina(n4630), .dinb(n4629), .dout(\result[59] ));
  jor  g3990(.dina(\address[1] ), .dinb(n3491), .dout(n4632));
  jor  g3991(.dina(n4452), .dinb(n3495), .dout(n4633));
  jand g3992(.dina(n4633), .dinb(n4632), .dout(\result[60] ));
  jor  g3993(.dina(\address[1] ), .dinb(n3448), .dout(n4635));
  jor  g3994(.dina(n4452), .dinb(n3452), .dout(n4636));
  jand g3995(.dina(n4636), .dinb(n4635), .dout(\result[61] ));
  jor  g3996(.dina(\address[1] ), .dinb(n3467), .dout(n4638));
  jor  g3997(.dina(n4452), .dinb(n3464), .dout(n4639));
  jand g3998(.dina(n4639), .dinb(n4638), .dout(\result[62] ));
  jor  g3999(.dina(\address[1] ), .dinb(n3456), .dout(n4641));
  jor  g4000(.dina(n4452), .dinb(n3460), .dout(n4642));
  jand g4001(.dina(n4642), .dinb(n4641), .dout(\result[63] ));
  jor  g4002(.dina(\address[1] ), .dinb(n3569), .dout(n4644));
  jor  g4003(.dina(n4452), .dinb(n3566), .dout(n4645));
  jand g4004(.dina(n4645), .dinb(n4644), .dout(\result[64] ));
  jor  g4005(.dina(\address[1] ), .dinb(n3558), .dout(n4647));
  jor  g4006(.dina(n4452), .dinb(n3562), .dout(n4648));
  jand g4007(.dina(n4648), .dinb(n4647), .dout(\result[65] ));
  jor  g4008(.dina(\address[1] ), .dinb(n3552), .dout(n4650));
  jor  g4009(.dina(n4452), .dinb(n3549), .dout(n4651));
  jand g4010(.dina(n4651), .dinb(n4650), .dout(\result[66] ));
  jor  g4011(.dina(\address[1] ), .dinb(n3541), .dout(n4653));
  jor  g4012(.dina(n4452), .dinb(n3545), .dout(n4654));
  jand g4013(.dina(n4654), .dinb(n4653), .dout(\result[67] ));
  jor  g4014(.dina(\address[1] ), .dinb(n3587), .dout(n4656));
  jor  g4015(.dina(n4452), .dinb(n3591), .dout(n4657));
  jand g4016(.dina(n4657), .dinb(n4656), .dout(\result[68] ));
  jor  g4017(.dina(\address[1] ), .dinb(n3595), .dout(n4659));
  jor  g4018(.dina(n4452), .dinb(n3599), .dout(n4660));
  jand g4019(.dina(n4660), .dinb(n4659), .dout(\result[69] ));
  jor  g4020(.dina(\address[1] ), .dinb(n3614), .dout(n4662));
  jor  g4021(.dina(n4452), .dinb(n3611), .dout(n4663));
  jand g4022(.dina(n4663), .dinb(n4662), .dout(\result[70] ));
  jor  g4023(.dina(\address[1] ), .dinb(n3603), .dout(n4665));
  jor  g4024(.dina(n4452), .dinb(n3607), .dout(n4666));
  jand g4025(.dina(n4666), .dinb(n4665), .dout(\result[71] ));
  jor  g4026(.dina(\address[1] ), .dinb(n3661), .dout(n4668));
  jor  g4027(.dina(n4452), .dinb(n3658), .dout(n4669));
  jand g4028(.dina(n4669), .dinb(n4668), .dout(\result[72] ));
  jor  g4029(.dina(\address[1] ), .dinb(n3650), .dout(n4671));
  jor  g4030(.dina(n4452), .dinb(n3654), .dout(n4672));
  jand g4031(.dina(n4672), .dinb(n4671), .dout(\result[73] ));
  jor  g4032(.dina(\address[1] ), .dinb(n3644), .dout(n4674));
  jor  g4033(.dina(n4452), .dinb(n3641), .dout(n4675));
  jand g4034(.dina(n4675), .dinb(n4674), .dout(\result[74] ));
  jor  g4035(.dina(\address[1] ), .dinb(n3633), .dout(n4677));
  jor  g4036(.dina(n4452), .dinb(n3637), .dout(n4678));
  jand g4037(.dina(n4678), .dinb(n4677), .dout(\result[75] ));
  jor  g4038(.dina(\address[1] ), .dinb(n3679), .dout(n4680));
  jor  g4039(.dina(n4452), .dinb(n3683), .dout(n4681));
  jand g4040(.dina(n4681), .dinb(n4680), .dout(\result[76] ));
  jor  g4041(.dina(\address[1] ), .dinb(n3687), .dout(n4683));
  jor  g4042(.dina(n4452), .dinb(n3691), .dout(n4684));
  jand g4043(.dina(n4684), .dinb(n4683), .dout(\result[77] ));
  jor  g4044(.dina(\address[1] ), .dinb(n3706), .dout(n4686));
  jor  g4045(.dina(n4452), .dinb(n3703), .dout(n4687));
  jand g4046(.dina(n4687), .dinb(n4686), .dout(\result[78] ));
  jor  g4047(.dina(\address[1] ), .dinb(n3695), .dout(n4689));
  jor  g4048(.dina(n4452), .dinb(n3699), .dout(n4690));
  jand g4049(.dina(n4690), .dinb(n4689), .dout(\result[79] ));
  jor  g4050(.dina(\address[1] ), .dinb(n3753), .dout(n4692));
  jor  g4051(.dina(n4452), .dinb(n3750), .dout(n4693));
  jand g4052(.dina(n4693), .dinb(n4692), .dout(\result[80] ));
  jor  g4053(.dina(\address[1] ), .dinb(n3742), .dout(n4695));
  jor  g4054(.dina(n4452), .dinb(n3746), .dout(n4696));
  jand g4055(.dina(n4696), .dinb(n4695), .dout(\result[81] ));
  jor  g4056(.dina(\address[1] ), .dinb(n3736), .dout(n4698));
  jor  g4057(.dina(n4452), .dinb(n3733), .dout(n4699));
  jand g4058(.dina(n4699), .dinb(n4698), .dout(\result[82] ));
  jor  g4059(.dina(\address[1] ), .dinb(n3725), .dout(n4701));
  jor  g4060(.dina(n4452), .dinb(n3729), .dout(n4702));
  jand g4061(.dina(n4702), .dinb(n4701), .dout(\result[83] ));
  jor  g4062(.dina(\address[1] ), .dinb(n3771), .dout(n4704));
  jor  g4063(.dina(n4452), .dinb(n3775), .dout(n4705));
  jand g4064(.dina(n4705), .dinb(n4704), .dout(\result[84] ));
  jor  g4065(.dina(\address[1] ), .dinb(n3779), .dout(n4707));
  jor  g4066(.dina(n4452), .dinb(n3783), .dout(n4708));
  jand g4067(.dina(n4708), .dinb(n4707), .dout(\result[85] ));
  jor  g4068(.dina(\address[1] ), .dinb(n3798), .dout(n4710));
  jor  g4069(.dina(n4452), .dinb(n3795), .dout(n4711));
  jand g4070(.dina(n4711), .dinb(n4710), .dout(\result[86] ));
  jor  g4071(.dina(\address[1] ), .dinb(n3787), .dout(n4713));
  jor  g4072(.dina(n4452), .dinb(n3791), .dout(n4714));
  jand g4073(.dina(n4714), .dinb(n4713), .dout(\result[87] ));
  jor  g4074(.dina(\address[1] ), .dinb(n3845), .dout(n4716));
  jor  g4075(.dina(n4452), .dinb(n3842), .dout(n4717));
  jand g4076(.dina(n4717), .dinb(n4716), .dout(\result[88] ));
  jor  g4077(.dina(\address[1] ), .dinb(n3834), .dout(n4719));
  jor  g4078(.dina(n4452), .dinb(n3838), .dout(n4720));
  jand g4079(.dina(n4720), .dinb(n4719), .dout(\result[89] ));
  jor  g4080(.dina(\address[1] ), .dinb(n3828), .dout(n4722));
  jor  g4081(.dina(n4452), .dinb(n3825), .dout(n4723));
  jand g4082(.dina(n4723), .dinb(n4722), .dout(\result[90] ));
  jor  g4083(.dina(\address[1] ), .dinb(n3817), .dout(n4725));
  jor  g4084(.dina(n4452), .dinb(n3821), .dout(n4726));
  jand g4085(.dina(n4726), .dinb(n4725), .dout(\result[91] ));
  jor  g4086(.dina(\address[1] ), .dinb(n3863), .dout(n4728));
  jor  g4087(.dina(n4452), .dinb(n3867), .dout(n4729));
  jand g4088(.dina(n4729), .dinb(n4728), .dout(\result[92] ));
  jor  g4089(.dina(\address[1] ), .dinb(n3871), .dout(n4731));
  jor  g4090(.dina(n4452), .dinb(n3875), .dout(n4732));
  jand g4091(.dina(n4732), .dinb(n4731), .dout(\result[93] ));
  jor  g4092(.dina(\address[1] ), .dinb(n3890), .dout(n4734));
  jor  g4093(.dina(n4452), .dinb(n3887), .dout(n4735));
  jand g4094(.dina(n4735), .dinb(n4734), .dout(\result[94] ));
  jor  g4095(.dina(\address[1] ), .dinb(n3879), .dout(n4737));
  jor  g4096(.dina(n4452), .dinb(n3883), .dout(n4738));
  jand g4097(.dina(n4738), .dinb(n4737), .dout(\result[95] ));
  jor  g4098(.dina(\address[1] ), .dinb(n3937), .dout(n4740));
  jor  g4099(.dina(n4452), .dinb(n3934), .dout(n4741));
  jand g4100(.dina(n4741), .dinb(n4740), .dout(\result[96] ));
  jor  g4101(.dina(\address[1] ), .dinb(n3926), .dout(n4743));
  jor  g4102(.dina(n4452), .dinb(n3930), .dout(n4744));
  jand g4103(.dina(n4744), .dinb(n4743), .dout(\result[97] ));
  jor  g4104(.dina(\address[1] ), .dinb(n3920), .dout(n4746));
  jor  g4105(.dina(n4452), .dinb(n3917), .dout(n4747));
  jand g4106(.dina(n4747), .dinb(n4746), .dout(\result[98] ));
  jor  g4107(.dina(\address[1] ), .dinb(n3909), .dout(n4749));
  jor  g4108(.dina(n4452), .dinb(n3913), .dout(n4750));
  jand g4109(.dina(n4750), .dinb(n4749), .dout(\result[99] ));
  jor  g4110(.dina(\address[1] ), .dinb(n3955), .dout(n4752));
  jor  g4111(.dina(n4452), .dinb(n3959), .dout(n4753));
  jand g4112(.dina(n4753), .dinb(n4752), .dout(\result[100] ));
  jor  g4113(.dina(\address[1] ), .dinb(n3963), .dout(n4755));
  jor  g4114(.dina(n4452), .dinb(n3967), .dout(n4756));
  jand g4115(.dina(n4756), .dinb(n4755), .dout(\result[101] ));
  jor  g4116(.dina(\address[1] ), .dinb(n3982), .dout(n4758));
  jor  g4117(.dina(n4452), .dinb(n3979), .dout(n4759));
  jand g4118(.dina(n4759), .dinb(n4758), .dout(\result[102] ));
  jor  g4119(.dina(\address[1] ), .dinb(n3971), .dout(n4761));
  jor  g4120(.dina(n4452), .dinb(n3975), .dout(n4762));
  jand g4121(.dina(n4762), .dinb(n4761), .dout(\result[103] ));
  jor  g4122(.dina(\address[1] ), .dinb(n4029), .dout(n4764));
  jor  g4123(.dina(n4452), .dinb(n4026), .dout(n4765));
  jand g4124(.dina(n4765), .dinb(n4764), .dout(\result[104] ));
  jor  g4125(.dina(\address[1] ), .dinb(n4018), .dout(n4767));
  jor  g4126(.dina(n4452), .dinb(n4022), .dout(n4768));
  jand g4127(.dina(n4768), .dinb(n4767), .dout(\result[105] ));
  jor  g4128(.dina(\address[1] ), .dinb(n4012), .dout(n4770));
  jor  g4129(.dina(n4452), .dinb(n4009), .dout(n4771));
  jand g4130(.dina(n4771), .dinb(n4770), .dout(\result[106] ));
  jor  g4131(.dina(\address[1] ), .dinb(n4001), .dout(n4773));
  jor  g4132(.dina(n4452), .dinb(n4005), .dout(n4774));
  jand g4133(.dina(n4774), .dinb(n4773), .dout(\result[107] ));
  jor  g4134(.dina(\address[1] ), .dinb(n4047), .dout(n4776));
  jor  g4135(.dina(n4452), .dinb(n4051), .dout(n4777));
  jand g4136(.dina(n4777), .dinb(n4776), .dout(\result[108] ));
  jor  g4137(.dina(\address[1] ), .dinb(n4055), .dout(n4779));
  jor  g4138(.dina(n4452), .dinb(n4059), .dout(n4780));
  jand g4139(.dina(n4780), .dinb(n4779), .dout(\result[109] ));
  jor  g4140(.dina(\address[1] ), .dinb(n4074), .dout(n4782));
  jor  g4141(.dina(n4452), .dinb(n4071), .dout(n4783));
  jand g4142(.dina(n4783), .dinb(n4782), .dout(\result[110] ));
  jor  g4143(.dina(\address[1] ), .dinb(n4063), .dout(n4785));
  jor  g4144(.dina(n4452), .dinb(n4067), .dout(n4786));
  jand g4145(.dina(n4786), .dinb(n4785), .dout(\result[111] ));
  jor  g4146(.dina(\address[1] ), .dinb(n4121), .dout(n4788));
  jor  g4147(.dina(n4452), .dinb(n4118), .dout(n4789));
  jand g4148(.dina(n4789), .dinb(n4788), .dout(\result[112] ));
  jor  g4149(.dina(\address[1] ), .dinb(n4110), .dout(n4791));
  jor  g4150(.dina(n4452), .dinb(n4114), .dout(n4792));
  jand g4151(.dina(n4792), .dinb(n4791), .dout(\result[113] ));
  jor  g4152(.dina(\address[1] ), .dinb(n4104), .dout(n4794));
  jor  g4153(.dina(n4452), .dinb(n4101), .dout(n4795));
  jand g4154(.dina(n4795), .dinb(n4794), .dout(\result[114] ));
  jor  g4155(.dina(\address[1] ), .dinb(n4093), .dout(n4797));
  jor  g4156(.dina(n4452), .dinb(n4097), .dout(n4798));
  jand g4157(.dina(n4798), .dinb(n4797), .dout(\result[115] ));
  jor  g4158(.dina(\address[1] ), .dinb(n4139), .dout(n4800));
  jor  g4159(.dina(n4452), .dinb(n4143), .dout(n4801));
  jand g4160(.dina(n4801), .dinb(n4800), .dout(\result[116] ));
  jor  g4161(.dina(\address[1] ), .dinb(n4147), .dout(n4803));
  jor  g4162(.dina(n4452), .dinb(n4151), .dout(n4804));
  jand g4163(.dina(n4804), .dinb(n4803), .dout(\result[117] ));
  jor  g4164(.dina(\address[1] ), .dinb(n4166), .dout(n4806));
  jor  g4165(.dina(n4452), .dinb(n4163), .dout(n4807));
  jand g4166(.dina(n4807), .dinb(n4806), .dout(\result[118] ));
  jor  g4167(.dina(\address[1] ), .dinb(n4155), .dout(n4809));
  jor  g4168(.dina(n4452), .dinb(n4159), .dout(n4810));
  jand g4169(.dina(n4810), .dinb(n4809), .dout(\result[119] ));
  jor  g4170(.dina(\address[1] ), .dinb(n4213), .dout(n4812));
  jor  g4171(.dina(n4452), .dinb(n4210), .dout(n4813));
  jand g4172(.dina(n4813), .dinb(n4812), .dout(\result[120] ));
  jor  g4173(.dina(\address[1] ), .dinb(n4202), .dout(n4815));
  jor  g4174(.dina(n4452), .dinb(n4206), .dout(n4816));
  jand g4175(.dina(n4816), .dinb(n4815), .dout(\result[121] ));
  jor  g4176(.dina(\address[1] ), .dinb(n4196), .dout(n4818));
  jor  g4177(.dina(n4452), .dinb(n4193), .dout(n4819));
  jand g4178(.dina(n4819), .dinb(n4818), .dout(\result[122] ));
  jor  g4179(.dina(\address[1] ), .dinb(n4185), .dout(n4821));
  jor  g4180(.dina(n4452), .dinb(n4189), .dout(n4822));
  jand g4181(.dina(n4822), .dinb(n4821), .dout(\result[123] ));
  jor  g4182(.dina(\address[1] ), .dinb(n4252), .dout(n4824));
  jor  g4183(.dina(n4452), .dinb(n4256), .dout(n4825));
  jand g4184(.dina(n4825), .dinb(n4824), .dout(\result[124] ));
  jor  g4185(.dina(\address[1] ), .dinb(n4239), .dout(n4827));
  jor  g4186(.dina(n4452), .dinb(n4243), .dout(n4828));
  jand g4187(.dina(n4828), .dinb(n4827), .dout(\result[125] ));
  jor  g4188(.dina(\address[1] ), .dinb(n4231), .dout(n4830));
  jor  g4189(.dina(n4452), .dinb(n4235), .dout(n4831));
  jand g4190(.dina(n4831), .dinb(n4830), .dout(\result[126] ));
  jand g4191(.dina(n4248), .dinb(n4246), .dout(\result[127] ));
  jor  g4192(.dina(\address[1] ), .dinb(n2783), .dout(n4834));
  jor  g4193(.dina(n4452), .dinb(n1711), .dout(n4835));
  jand g4194(.dina(n4835), .dinb(n4834), .dout(\address[0] ));
endmodule


