/*

c499:
	jxor: 108
	jspl: 34
	jspl3: 68
	jnot: 17
	jcb: 10
	jdff: 382
	jand: 61

Summary:
	jxor: 108
	jspl: 34
	jspl3: 68
	jnot: 17
	jcb: 10
	jdff: 382
	jand: 61
*/

module c499(gclk, Gid0, Gid1, Gid2, Gid3, Gid4, Gid5, Gid6, Gid7, Gid8, Gid9, Gid10, Gid11, Gid12, Gid13, Gid14, Gid15, Gid16, Gid17, Gid18, Gid19, Gid20, Gid21, Gid22, Gid23, Gid24, Gid25, Gid26, Gid27, Gid28, Gid29, Gid30, Gid31, Gic0, Gic1, Gic2, Gic3, Gic4, Gic5, Gic6, Gic7, Gr, God0, God1, God2, God3, God4, God5, God6, God7, God8, God9, God10, God11, God12, God13, God14, God15, God16, God17, God18, God19, God20, God21, God22, God23, God24, God25, God26, God27, God28, God29, God30, God31);
	input gclk;
	input Gid0;
	input Gid1;
	input Gid2;
	input Gid3;
	input Gid4;
	input Gid5;
	input Gid6;
	input Gid7;
	input Gid8;
	input Gid9;
	input Gid10;
	input Gid11;
	input Gid12;
	input Gid13;
	input Gid14;
	input Gid15;
	input Gid16;
	input Gid17;
	input Gid18;
	input Gid19;
	input Gid20;
	input Gid21;
	input Gid22;
	input Gid23;
	input Gid24;
	input Gid25;
	input Gid26;
	input Gid27;
	input Gid28;
	input Gid29;
	input Gid30;
	input Gid31;
	input Gic0;
	input Gic1;
	input Gic2;
	input Gic3;
	input Gic4;
	input Gic5;
	input Gic6;
	input Gic7;
	input Gr;
	output God0;
	output God1;
	output God2;
	output God3;
	output God4;
	output God5;
	output God6;
	output God7;
	output God8;
	output God9;
	output God10;
	output God11;
	output God12;
	output God13;
	output God14;
	output God15;
	output God16;
	output God17;
	output God18;
	output God19;
	output God20;
	output God21;
	output God22;
	output God23;
	output God24;
	output God25;
	output God26;
	output God27;
	output God28;
	output God29;
	output God30;
	output God31;
	wire n73;
	wire n74;
	wire n75;
	wire n76;
	wire n77;
	wire n78;
	wire n79;
	wire n80;
	wire n81;
	wire n82;
	wire n83;
	wire n84;
	wire n85;
	wire n86;
	wire n87;
	wire n88;
	wire n89;
	wire n90;
	wire n91;
	wire n92;
	wire n93;
	wire n94;
	wire n95;
	wire n96;
	wire n97;
	wire n98;
	wire n99;
	wire n100;
	wire n101;
	wire n102;
	wire n103;
	wire n104;
	wire n105;
	wire n106;
	wire n107;
	wire n108;
	wire n109;
	wire n110;
	wire n111;
	wire n112;
	wire n113;
	wire n114;
	wire n115;
	wire n116;
	wire n117;
	wire n118;
	wire n119;
	wire n120;
	wire n121;
	wire n122;
	wire n123;
	wire n124;
	wire n125;
	wire n126;
	wire n127;
	wire n128;
	wire n129;
	wire n130;
	wire n131;
	wire n132;
	wire n133;
	wire n134;
	wire n135;
	wire n136;
	wire n137;
	wire n138;
	wire n139;
	wire n140;
	wire n141;
	wire n142;
	wire n143;
	wire n144;
	wire n145;
	wire n146;
	wire n147;
	wire n148;
	wire n149;
	wire n150;
	wire n151;
	wire n152;
	wire n153;
	wire n154;
	wire n155;
	wire n156;
	wire n157;
	wire n158;
	wire n159;
	wire n160;
	wire n161;
	wire n162;
	wire n163;
	wire n164;
	wire n165;
	wire n166;
	wire n167;
	wire n168;
	wire n169;
	wire n170;
	wire n171;
	wire n172;
	wire n173;
	wire n174;
	wire n175;
	wire n176;
	wire n178;
	wire n179;
	wire n181;
	wire n182;
	wire n184;
	wire n185;
	wire n187;
	wire n188;
	wire n189;
	wire n190;
	wire n192;
	wire n194;
	wire n196;
	wire n198;
	wire n199;
	wire n200;
	wire n201;
	wire n202;
	wire n204;
	wire n206;
	wire n208;
	wire n210;
	wire n211;
	wire n212;
	wire n214;
	wire n216;
	wire n218;
	wire n220;
	wire n221;
	wire n222;
	wire n223;
	wire n224;
	wire n225;
	wire n226;
	wire n227;
	wire n228;
	wire n229;
	wire n230;
	wire n231;
	wire n233;
	wire n235;
	wire n237;
	wire n239;
	wire n240;
	wire n241;
	wire n242;
	wire n244;
	wire n246;
	wire n248;
	wire n250;
	wire n251;
	wire n252;
	wire n254;
	wire n256;
	wire n258;
	wire n260;
	wire n261;
	wire n263;
	wire n265;
	wire n267;
	wire [2:0] w_Gid0_0;
	wire [2:0] w_Gid1_0;
	wire [2:0] w_Gid2_0;
	wire [2:0] w_Gid3_0;
	wire [2:0] w_Gid4_0;
	wire [2:0] w_Gid5_0;
	wire [2:0] w_Gid6_0;
	wire [2:0] w_Gid7_0;
	wire [2:0] w_Gid8_0;
	wire [2:0] w_Gid9_0;
	wire [2:0] w_Gid10_0;
	wire [2:0] w_Gid11_0;
	wire [2:0] w_Gid12_0;
	wire [2:0] w_Gid13_0;
	wire [2:0] w_Gid14_0;
	wire [2:0] w_Gid15_0;
	wire [2:0] w_Gid16_0;
	wire [2:0] w_Gid17_0;
	wire [2:0] w_Gid18_0;
	wire [2:0] w_Gid19_0;
	wire [2:0] w_Gid20_0;
	wire [2:0] w_Gid21_0;
	wire [2:0] w_Gid22_0;
	wire [2:0] w_Gid23_0;
	wire [2:0] w_Gid24_0;
	wire [2:0] w_Gid25_0;
	wire [2:0] w_Gid26_0;
	wire [2:0] w_Gid27_0;
	wire [2:0] w_Gid28_0;
	wire [2:0] w_Gid29_0;
	wire [2:0] w_Gid30_0;
	wire [2:0] w_Gid31_0;
	wire [2:0] w_n74_0;
	wire [2:0] w_n74_1;
	wire [2:0] w_n74_2;
	wire [1:0] w_n74_3;
	wire [1:0] w_n78_0;
	wire [1:0] w_n85_0;
	wire [2:0] w_n87_0;
	wire [1:0] w_n87_1;
	wire [2:0] w_n88_0;
	wire [2:0] w_n88_1;
	wire [1:0] w_n93_0;
	wire [1:0] w_n97_0;
	wire [2:0] w_n102_0;
	wire [1:0] w_n102_1;
	wire [1:0] w_n107_0;
	wire [1:0] w_n111_0;
	wire [2:0] w_n116_0;
	wire [1:0] w_n116_1;
	wire [2:0] w_n117_0;
	wire [2:0] w_n117_1;
	wire [1:0] w_n118_0;
	wire [2:0] w_n126_0;
	wire [1:0] w_n126_1;
	wire [2:0] w_n127_0;
	wire [2:0] w_n127_1;
	wire [2:0] w_n135_0;
	wire [1:0] w_n135_1;
	wire [1:0] w_n141_0;
	wire [1:0] w_n145_0;
	wire [2:0] w_n150_0;
	wire [1:0] w_n150_1;
	wire [2:0] w_n159_0;
	wire [1:0] w_n159_1;
	wire [2:0] w_n167_0;
	wire [1:0] w_n167_1;
	wire [2:0] w_n173_0;
	wire [1:0] w_n174_0;
	wire [2:0] w_n175_0;
	wire [1:0] w_n175_1;
	wire [2:0] w_n178_0;
	wire [2:0] w_n178_1;
	wire [2:0] w_n181_0;
	wire [2:0] w_n181_1;
	wire [2:0] w_n184_0;
	wire [2:0] w_n184_1;
	wire [2:0] w_n187_0;
	wire [2:0] w_n187_1;
	wire [1:0] w_n188_0;
	wire [2:0] w_n189_0;
	wire [1:0] w_n189_1;
	wire [2:0] w_n198_0;
	wire [2:0] w_n198_1;
	wire [1:0] w_n199_0;
	wire [2:0] w_n201_0;
	wire [1:0] w_n201_1;
	wire [2:0] w_n211_0;
	wire [1:0] w_n211_1;
	wire [1:0] w_n220_0;
	wire [1:0] w_n228_0;
	wire [1:0] w_n229_0;
	wire [2:0] w_n230_0;
	wire [1:0] w_n230_1;
	wire [1:0] w_n240_0;
	wire [2:0] w_n241_0;
	wire [1:0] w_n241_1;
	wire [1:0] w_n250_0;
	wire [2:0] w_n251_0;
	wire [1:0] w_n251_1;
	wire [2:0] w_n260_0;
	wire [1:0] w_n260_1;
	wire w_dff_A_Gay8MZ4x5_1;
	wire w_dff_A_8UoaUcmQ7_1;
	wire w_dff_A_nkkr6ssB2_0;
	wire w_dff_A_SoPSj0JI0_1;
	wire w_dff_A_z8wTnRGS4_0;
	wire w_dff_A_p0OCm6EC3_0;
	wire w_dff_A_iUsVz9Of4_0;
	wire w_dff_A_D2t15BiB9_1;
	wire w_dff_A_VvqVNZHs2_1;
	wire w_dff_A_AFC26J8h4_1;
	wire w_dff_A_gL4MMgIh2_0;
	wire w_dff_A_VflmckS26_0;
	wire w_dff_A_obfMM42W9_0;
	wire w_dff_A_WxCg7RGe8_1;
	wire w_dff_A_dVq2s78T0_1;
	wire w_dff_A_ybqClvk39_1;
	wire w_dff_A_mlZA7mzT3_0;
	wire w_dff_A_m3AhxUKP9_0;
	wire w_dff_A_RdyzR5Yi3_0;
	wire w_dff_A_lfU4Xgec4_1;
	wire w_dff_A_E0PG8tGi1_1;
	wire w_dff_A_k5aMHF8R6_1;
	wire w_dff_B_ZNirXdbH6_2;
	wire w_dff_A_j4XMoKDy1_0;
	wire w_dff_A_gfYr5qa00_0;
	wire w_dff_A_7HOZnrRL8_0;
	wire w_dff_A_a0CkAKZ58_2;
	wire w_dff_A_we2xVxLm6_2;
	wire w_dff_A_cMWeQ5XI8_2;
	wire w_dff_A_zKjvttGZ3_0;
	wire w_dff_A_xNDejBvk0_0;
	wire w_dff_A_WAcsnX4T5_0;
	wire w_dff_A_MLKUktyu2_1;
	wire w_dff_A_mZ7wmJHc4_1;
	wire w_dff_A_cru1nvzF8_1;
	wire w_dff_A_t8diCatx3_0;
	wire w_dff_A_FEisqJMX8_0;
	wire w_dff_A_TSdGAzNV8_0;
	wire w_dff_A_MAsuxIbO7_2;
	wire w_dff_A_3T3QLBvE1_2;
	wire w_dff_A_JArBfUQ79_2;
	wire w_dff_A_vio35cWh5_1;
	wire w_dff_A_36jn2a659_1;
	wire w_dff_A_QP3bYQP69_1;
	wire w_dff_A_g3WR95nz3_2;
	wire w_dff_A_jkOEhk0c1_2;
	wire w_dff_A_jozhULJA9_2;
	wire w_dff_A_6fvZ8SAh2_0;
	wire w_dff_A_GQdN42S37_1;
	wire w_dff_A_FOg1v7fp9_1;
	wire w_dff_A_wxGtXfff4_1;
	wire w_dff_A_iJoDg3Ir3_2;
	wire w_dff_A_C72QquDl7_2;
	wire w_dff_A_I8uXnHgx3_2;
	wire w_dff_A_o7MXsCVg9_1;
	wire w_dff_A_ohslviSy4_1;
	wire w_dff_A_uB2Dc9v70_1;
	wire w_dff_A_VJiCPsNs4_1;
	wire w_dff_A_ONG3ilCy9_2;
	wire w_dff_A_bmfCiTBG4_2;
	wire w_dff_A_umK8VC3f9_2;
	wire w_dff_A_QG81S6Au8_0;
	wire w_dff_B_ubnJPw2i5_0;
	wire w_dff_B_nYQA3b499_0;
	wire w_dff_B_qL0lohj90_1;
	wire w_dff_A_ZwEhqkxI7_1;
	wire w_dff_A_4NXxozkh3_0;
	wire w_dff_A_Lr87YYC90_0;
	wire w_dff_A_8yOhhC1f0_0;
	wire w_dff_A_M1h9aFMj4_0;
	wire w_dff_A_i9j5lDzb9_0;
	wire w_dff_A_vGfJnd7g9_0;
	wire w_dff_A_do0Lp34X4_0;
	wire w_dff_A_bqk6m5BF1_0;
	wire w_dff_A_J2bJJcFI8_0;
	wire w_dff_A_Y7lcpacD6_0;
	wire w_dff_A_hhVzoZaR9_0;
	wire w_dff_A_P6cRG2mZ2_0;
	wire w_dff_A_EMu4TDRX3_0;
	wire w_dff_A_AK3xpoD71_0;
	wire w_dff_A_xFjWKTk92_0;
	wire w_dff_A_paJVS0G39_0;
	wire w_dff_A_8VO8diVD1_0;
	wire w_dff_A_asTtwopN9_0;
	wire w_dff_B_i2Mv9mSE2_0;
	wire w_dff_A_7unGc1N81_0;
	wire w_dff_A_Ift1tEiP2_0;
	wire w_dff_A_WhzBcMHk9_0;
	wire w_dff_A_QRlEQHcp2_2;
	wire w_dff_A_fGHsChWy1_2;
	wire w_dff_A_F0a4qMEL1_2;
	wire w_dff_A_USYzVecP0_1;
	wire w_dff_A_rIbjrGUp0_0;
	wire w_dff_A_FMIl07QG2_0;
	wire w_dff_A_9OeaZVPh4_0;
	wire w_dff_A_jUt0qhEZ6_0;
	wire w_dff_A_HWifq8Fu0_0;
	wire w_dff_A_O0Z7EDWG0_0;
	wire w_dff_A_9WsiYxJS2_0;
	wire w_dff_A_3y2Q2Tqr1_0;
	wire w_dff_A_Lni5NrPW5_0;
	wire w_dff_A_cYKSY5fp6_0;
	wire w_dff_A_ZkJbhuKU3_0;
	wire w_dff_A_dRNxF2B02_0;
	wire w_dff_A_k5Rv8Bkw2_0;
	wire w_dff_A_kjRatyLr2_0;
	wire w_dff_A_o23deXt75_0;
	wire w_dff_A_L1GO89uh6_0;
	wire w_dff_A_srLF8pSZ3_0;
	wire w_dff_A_jJuM7kdD5_0;
	wire w_dff_B_nOPe9sMB7_0;
	wire w_dff_B_UC88yyfr6_2;
	wire w_dff_A_7GG0Pdeh6_0;
	wire w_dff_A_W1UZUwC65_0;
	wire w_dff_A_d3Pa53nW2_0;
	wire w_dff_A_AaNgmwLP3_2;
	wire w_dff_A_8iiCmORe1_2;
	wire w_dff_A_vdMCMSdo5_2;
	wire w_dff_A_7VTeUlZZ6_1;
	wire w_dff_A_eIv5XzI46_0;
	wire w_dff_A_O76DOFuz5_0;
	wire w_dff_A_A4go7Xc77_0;
	wire w_dff_A_6NZCI8ZK6_0;
	wire w_dff_A_j2adSQB68_0;
	wire w_dff_A_djVnZcu11_0;
	wire w_dff_A_Ug0wiIoZ7_0;
	wire w_dff_A_3lXIVw5j2_0;
	wire w_dff_A_KnxHH5LI4_0;
	wire w_dff_A_1dR3VcGE8_0;
	wire w_dff_A_PLZhoxte0_0;
	wire w_dff_A_tlO5yp5z1_0;
	wire w_dff_A_gSm9D3Ag9_0;
	wire w_dff_A_Sq4JzbZU8_0;
	wire w_dff_A_V7qKu6Bj9_0;
	wire w_dff_A_PyxwTlgq3_0;
	wire w_dff_A_eZFHzSBZ1_0;
	wire w_dff_A_ibDwxNCx3_0;
	wire w_dff_A_lxrLuyYV2_0;
	wire w_dff_A_HaVaPBOT7_0;
	wire w_dff_A_MbULmuV91_0;
	wire w_dff_A_FCbjU2kj8_0;
	wire w_dff_A_y728LCBF3_0;
	wire w_dff_A_wRXh8FI02_0;
	wire w_dff_A_4tyfHfTH3_0;
	wire w_dff_A_RflG3I773_0;
	wire w_dff_A_mLEMYJRM9_0;
	wire w_dff_A_MRxFezn76_0;
	wire w_dff_A_AnF5QnyT9_0;
	wire w_dff_A_pxK0fo0l9_0;
	wire w_dff_A_slVlHIJ22_0;
	wire w_dff_A_UhdG2aDJ3_0;
	wire w_dff_A_qf8HLpB87_0;
	wire w_dff_A_hk1hBb262_0;
	wire w_dff_A_s3aYkSp83_0;
	wire w_dff_A_p0JsYRz87_0;
	wire w_dff_A_lD0vxeIb6_0;
	wire w_dff_A_zVPlDPcz1_0;
	wire w_dff_A_Szl2p8Dp3_0;
	wire w_dff_A_y2fbIcPa9_0;
	wire w_dff_A_ZIWQSUWm1_0;
	wire w_dff_A_0mxIEL0Z9_0;
	wire w_dff_A_ZeTrkn1Q2_0;
	wire w_dff_A_kdFYze5e1_0;
	wire w_dff_A_2bZYM1jj9_0;
	wire w_dff_B_fq2pqfIy1_1;
	wire w_dff_A_PrT5yRJK7_0;
	wire w_dff_A_K4S6b3Qc3_0;
	wire w_dff_A_oPbRgCbe7_0;
	wire w_dff_A_6k88Ow9F8_0;
	wire w_dff_A_JJJrjD4X6_0;
	wire w_dff_A_4iWHi9c62_0;
	wire w_dff_A_JmYSlVj16_0;
	wire w_dff_A_9f7E5E7Q2_0;
	wire w_dff_A_PGuNR5kM5_0;
	wire w_dff_A_Ks24DUMm1_0;
	wire w_dff_A_2b1dVPwE6_0;
	wire w_dff_A_OR7hYgjl6_0;
	wire w_dff_A_dn89tSFB9_0;
	wire w_dff_A_A0n2jZf65_0;
	wire w_dff_A_EqzUeRIk8_0;
	wire w_dff_A_Uj4GsI588_0;
	wire w_dff_A_LWVePi6g3_0;
	wire w_dff_A_lpdSTX472_0;
	wire w_dff_A_x2JCpfEA2_0;
	wire w_dff_A_CRzMu6Ej3_0;
	wire w_dff_A_t0ciBwgo1_0;
	wire w_dff_A_HgWc9BkZ2_0;
	wire w_dff_A_KIJqRfKM4_0;
	wire w_dff_A_2vN6qVH66_0;
	wire w_dff_A_tavcwFC29_0;
	wire w_dff_A_ALXC0HG02_0;
	wire w_dff_A_KqvraJus8_0;
	wire w_dff_A_PXTVRGeM9_1;
	wire w_dff_A_1FxENjWr2_0;
	wire w_dff_A_ogf2vX5S4_0;
	wire w_dff_A_jqihCHYU0_0;
	wire w_dff_A_T0SHlAxV4_0;
	wire w_dff_A_WFMAe56z7_0;
	wire w_dff_A_kTa85LaC5_0;
	wire w_dff_A_uvTLUANg3_0;
	wire w_dff_A_gZbEjkNZ1_0;
	wire w_dff_A_ZlF6DRNS8_0;
	wire w_dff_A_tiBLV1YL1_0;
	wire w_dff_A_1rqcKS623_0;
	wire w_dff_A_FovqzTDo5_0;
	wire w_dff_A_ObNp9zp69_0;
	wire w_dff_A_YJG9NDrE3_0;
	wire w_dff_A_Zwo4CKf33_0;
	wire w_dff_A_rx7JAJlH8_0;
	wire w_dff_A_nhJEgkeJ4_0;
	wire w_dff_A_SBxBORC27_0;
	wire w_dff_A_tV8yo2h87_0;
	wire w_dff_A_buwdRfLs2_0;
	wire w_dff_A_B0zqrSuL5_0;
	wire w_dff_A_eiyFXXyB3_0;
	wire w_dff_A_AggnXpA57_0;
	wire w_dff_A_t9LVRxAo2_0;
	wire w_dff_A_EhC0h2vs5_0;
	wire w_dff_A_j0D5SOUx4_0;
	wire w_dff_A_8AF4rwWG4_0;
	wire w_dff_A_0IZLWlvP1_0;
	wire w_dff_A_B860Ugzw7_0;
	wire w_dff_A_zgh7f9YY9_0;
	wire w_dff_A_GoHujcHd9_0;
	wire w_dff_A_GoZClivP6_0;
	wire w_dff_A_S8VSJANp4_0;
	wire w_dff_A_6YWNRBmi0_0;
	wire w_dff_A_Mo7Czp4I5_0;
	wire w_dff_A_Fm81bVXb4_0;
	wire w_dff_A_rTsSmuLl0_0;
	wire w_dff_A_5BQ3PXpO5_0;
	wire w_dff_A_WTIBzFbc1_0;
	wire w_dff_A_0JzMntPC8_0;
	wire w_dff_A_NogwJga58_0;
	wire w_dff_A_6pFiOnxD8_0;
	wire w_dff_A_eMP34gdl6_0;
	wire w_dff_A_vFmJqvz96_0;
	wire w_dff_A_jeIqdny36_0;
	wire w_dff_B_cIPsQN239_1;
	wire w_dff_A_LWCSZxky9_0;
	wire w_dff_A_CtBCDOTn2_0;
	wire w_dff_A_0AKNiRU74_0;
	wire w_dff_A_r4oiOSDq0_0;
	wire w_dff_A_YDvw6Okc5_0;
	wire w_dff_A_yjVHrI783_0;
	wire w_dff_A_8aYyWgMp2_0;
	wire w_dff_A_hyVhuwv11_0;
	wire w_dff_A_pEGxduJo7_0;
	wire w_dff_A_YtPkck9X0_0;
	wire w_dff_A_3GW6Q84W5_0;
	wire w_dff_A_xlCckJXS9_0;
	wire w_dff_A_Eqxn9ihg9_0;
	wire w_dff_A_09sQ4T991_0;
	wire w_dff_A_jinmfTAn7_0;
	wire w_dff_A_tIx9bA3Q0_0;
	wire w_dff_A_w8A5x5PP4_0;
	wire w_dff_A_TLDVzjjS5_0;
	wire w_dff_A_Pm24qRSh2_0;
	wire w_dff_A_UQ6moDOL1_0;
	wire w_dff_A_DunxYemY2_0;
	wire w_dff_A_2aI3FGae6_0;
	wire w_dff_A_IsXqFmFF4_0;
	wire w_dff_A_561XGa8Q4_0;
	wire w_dff_A_XfgkVAcc8_0;
	wire w_dff_A_c6GpQIdt8_0;
	wire w_dff_A_7a90pXgD9_0;
	wire w_dff_A_k0bCiLaS2_1;
	wire w_dff_A_f2s8mWow7_1;
	wire w_dff_A_5g65sS2q0_1;
	wire w_dff_A_kCJ787kt9_2;
	wire w_dff_A_8aSTICIo0_2;
	wire w_dff_A_SI7LRVvI5_2;
	wire w_dff_A_onFBGz5h5_1;
	wire w_dff_A_ahfjs8qw3_0;
	wire w_dff_A_4CBE20Fx6_0;
	wire w_dff_A_CmfBq9W25_0;
	wire w_dff_A_VkDfYNUq3_0;
	wire w_dff_A_986HQcMu7_0;
	wire w_dff_A_7atJrpkP6_0;
	wire w_dff_A_wIzZywLv4_0;
	wire w_dff_A_2n5YP8lt9_0;
	wire w_dff_A_Mk7fOtus9_0;
	wire w_dff_A_Iobxln0X2_0;
	wire w_dff_A_y74magwy5_0;
	wire w_dff_A_EBxyZdkC6_0;
	wire w_dff_A_4WUkd2ps2_0;
	wire w_dff_A_glBX3B5F6_0;
	wire w_dff_A_aYEnnFAd7_0;
	wire w_dff_A_k6sA7Hxe1_0;
	wire w_dff_A_yhkskwpx8_0;
	wire w_dff_A_atPkpVhr5_0;
	wire w_dff_A_xQ0AQxpe6_0;
	wire w_dff_A_9X4gwM5a4_0;
	wire w_dff_A_lo9aW5vm6_0;
	wire w_dff_A_IVsM3AX00_0;
	wire w_dff_A_7WgGb0fo2_0;
	wire w_dff_A_v6WQ1kX65_0;
	wire w_dff_A_NDLb4voV1_0;
	wire w_dff_A_pXkblSMP7_0;
	wire w_dff_A_PiQJmDTh0_0;
	wire w_dff_A_Q4CMYELA8_0;
	wire w_dff_A_3YawHl5y3_0;
	wire w_dff_A_OKVBf5Ep3_0;
	wire w_dff_A_vqbeihJG0_0;
	wire w_dff_A_7rrmaD3S8_0;
	wire w_dff_A_aSyoe34x4_0;
	wire w_dff_A_ooiB0p4j7_0;
	wire w_dff_A_z4c8E6dp7_0;
	wire w_dff_A_nCnJAGQY6_0;
	wire w_dff_A_XpIpBYFo4_0;
	wire w_dff_A_SjxrMhjv6_0;
	wire w_dff_A_diQhLNkK8_0;
	wire w_dff_A_vLDnubxj3_0;
	wire w_dff_A_DNmO7cE60_0;
	wire w_dff_A_lXkyjtLR9_0;
	wire w_dff_A_dOzgrWnE1_0;
	wire w_dff_A_0eJjrkoH9_0;
	wire w_dff_A_4KrvNnKl3_0;
	wire w_dff_A_6wLaNSOi9_0;
	wire w_dff_A_2kyX6NGj2_0;
	wire w_dff_A_tGScyidT4_0;
	wire w_dff_A_fSged4Wv5_0;
	wire w_dff_A_Zi3qTDkl0_0;
	wire w_dff_A_QurSle926_0;
	wire w_dff_A_3LAcBKPj4_0;
	wire w_dff_A_4GZxTSrF7_0;
	wire w_dff_A_QIjOxqaN9_0;
	wire w_dff_A_vh1jU26g1_0;
	wire w_dff_A_q1lzO1Xl8_0;
	wire w_dff_A_MEyKYcYZ2_0;
	wire w_dff_A_GSX6na7u8_0;
	wire w_dff_A_2o412wT18_0;
	wire w_dff_A_C9yWhCjS6_0;
	wire w_dff_A_BeOAonQr0_0;
	wire w_dff_A_Vhb6DImv1_0;
	wire w_dff_A_iv4e9N5q4_0;
	wire w_dff_A_vjSqQ4gs1_0;
	wire w_dff_A_JuDPkQfu1_0;
	wire w_dff_A_Qv375HHq5_0;
	wire w_dff_A_QIqiZhg58_0;
	wire w_dff_A_BvHJu2zl3_0;
	wire w_dff_A_Asr8THu82_0;
	wire w_dff_A_oOqD5JSR8_0;
	wire w_dff_A_6pNqEd4X3_0;
	wire w_dff_A_1YGnxI0q7_0;
	wire w_dff_B_R4HEtQGW7_1;
	wire w_dff_A_OTrU2NfY0_0;
	wire w_dff_A_I9IxrMYY2_0;
	wire w_dff_A_4ojeLkYG9_0;
	wire w_dff_A_THSwPUtt4_0;
	wire w_dff_A_n2MoqrZ97_0;
	wire w_dff_A_l4Qsk1qB5_0;
	wire w_dff_A_i4dMAA0L4_0;
	wire w_dff_A_yMN71vaN3_0;
	wire w_dff_A_DMwycXsd8_0;
	wire w_dff_A_94bBd39p7_0;
	wire w_dff_A_hZhPAOVA3_0;
	wire w_dff_A_04XiGpaa8_0;
	wire w_dff_A_AJHbVk5w4_0;
	wire w_dff_A_hZcE0wOS9_0;
	wire w_dff_A_aOfOJiTD2_0;
	wire w_dff_A_OPBRgcvV5_0;
	wire w_dff_A_L0J8lgij4_0;
	wire w_dff_A_7fxMyzXe9_0;
	wire w_dff_A_caidO8Up4_0;
	wire w_dff_A_YY7WWgQg2_0;
	wire w_dff_A_5FUYyccq4_0;
	wire w_dff_A_CMouldip0_0;
	wire w_dff_A_XmXmT7pS5_0;
	wire w_dff_A_LqB4KDHE2_0;
	wire w_dff_A_tngNbI3j8_0;
	wire w_dff_A_JEOsdz1W0_0;
	wire w_dff_A_f4JIbIaN0_0;
	wire w_dff_A_BhjqQ1Cs2_0;
	wire w_dff_A_l71KpzS20_0;
	wire w_dff_A_VUtDisqQ5_0;
	wire w_dff_A_WaxHf69c0_0;
	wire w_dff_A_OiVHDl0Z6_0;
	wire w_dff_A_Z7zZaQM37_0;
	wire w_dff_A_HO71wEew0_0;
	wire w_dff_A_XRH2tvWv2_0;
	wire w_dff_A_D8w0sMRT0_0;
	jnot g000(.din(Gic0),.dout(n73),.clk(gclk));
	jnot g001(.din(Gr),.dout(n74),.clk(gclk));
	jcb g002(.dina(w_n74_3[1]),.dinb(n73),.dout(n75));
	jxor g003(.dina(w_Gid17_0[2]),.dinb(w_Gid16_0[2]),.dout(n76),.clk(gclk));
	jxor g004(.dina(w_Gid19_0[2]),.dinb(w_Gid18_0[2]),.dout(n77),.clk(gclk));
	jxor g005(.dina(n77),.dinb(n76),.dout(n78),.clk(gclk));
	jxor g006(.dina(w_n78_0[1]),.dinb(w_dff_B_cIPsQN239_1),.dout(n79),.clk(gclk));
	jxor g007(.dina(w_Gid4_0[2]),.dinb(w_Gid0_0[2]),.dout(n80),.clk(gclk));
	jxor g008(.dina(w_Gid12_0[2]),.dinb(w_Gid8_0[2]),.dout(n81),.clk(gclk));
	jxor g009(.dina(n81),.dinb(n80),.dout(n82),.clk(gclk));
	jxor g010(.dina(w_Gid21_0[2]),.dinb(w_Gid20_0[2]),.dout(n83),.clk(gclk));
	jxor g011(.dina(w_Gid23_0[2]),.dinb(w_Gid22_0[2]),.dout(n84),.clk(gclk));
	jxor g012(.dina(n84),.dinb(n83),.dout(n85),.clk(gclk));
	jxor g013(.dina(w_n85_0[1]),.dinb(n82),.dout(n86),.clk(gclk));
	jxor g014(.dina(n86),.dinb(n79),.dout(n87),.clk(gclk));
	jnot g015(.din(w_n87_1[1]),.dout(n88),.clk(gclk));
	jnot g016(.din(Gic7),.dout(n89),.clk(gclk));
	jcb g017(.dina(w_n74_3[0]),.dinb(n89),.dout(n90));
	jxor g018(.dina(w_Gid5_0[2]),.dinb(w_Gid4_0[1]),.dout(n91),.clk(gclk));
	jxor g019(.dina(w_Gid7_0[2]),.dinb(w_Gid6_0[2]),.dout(n92),.clk(gclk));
	jxor g020(.dina(n92),.dinb(n91),.dout(n93),.clk(gclk));
	jxor g021(.dina(w_n93_0[1]),.dinb(w_dff_B_R4HEtQGW7_1),.dout(n94),.clk(gclk));
	jxor g022(.dina(w_Gid13_0[2]),.dinb(w_Gid12_0[1]),.dout(n95),.clk(gclk));
	jxor g023(.dina(w_Gid15_0[2]),.dinb(w_Gid14_0[2]),.dout(n96),.clk(gclk));
	jxor g024(.dina(n96),.dinb(n95),.dout(n97),.clk(gclk));
	jxor g025(.dina(w_Gid23_0[1]),.dinb(w_Gid19_0[1]),.dout(n98),.clk(gclk));
	jxor g026(.dina(w_Gid31_0[2]),.dinb(w_Gid27_0[2]),.dout(n99),.clk(gclk));
	jxor g027(.dina(n99),.dinb(n98),.dout(n100),.clk(gclk));
	jxor g028(.dina(n100),.dinb(w_n97_0[1]),.dout(n101),.clk(gclk));
	jxor g029(.dina(n101),.dinb(n94),.dout(n102),.clk(gclk));
	jnot g030(.din(Gic6),.dout(n103),.clk(gclk));
	jcb g031(.dina(w_n74_2[2]),.dinb(n103),.dout(n104));
	jxor g032(.dina(w_Gid1_0[2]),.dinb(w_Gid0_0[1]),.dout(n105),.clk(gclk));
	jxor g033(.dina(w_Gid3_0[2]),.dinb(w_Gid2_0[2]),.dout(n106),.clk(gclk));
	jxor g034(.dina(n106),.dinb(n105),.dout(n107),.clk(gclk));
	jxor g035(.dina(w_n107_0[1]),.dinb(w_dff_B_qL0lohj90_1),.dout(n108),.clk(gclk));
	jxor g036(.dina(w_Gid9_0[2]),.dinb(w_Gid8_0[1]),.dout(n109),.clk(gclk));
	jxor g037(.dina(w_Gid11_0[2]),.dinb(w_Gid10_0[2]),.dout(n110),.clk(gclk));
	jxor g038(.dina(n110),.dinb(n109),.dout(n111),.clk(gclk));
	jxor g039(.dina(w_Gid22_0[1]),.dinb(w_Gid18_0[1]),.dout(n112),.clk(gclk));
	jxor g040(.dina(w_Gid30_0[2]),.dinb(w_Gid26_0[2]),.dout(n113),.clk(gclk));
	jxor g041(.dina(n113),.dinb(n112),.dout(n114),.clk(gclk));
	jxor g042(.dina(n114),.dinb(w_n111_0[1]),.dout(n115),.clk(gclk));
	jxor g043(.dina(n115),.dinb(n108),.dout(n116),.clk(gclk));
	jnot g044(.din(w_n116_1[1]),.dout(n117),.clk(gclk));
	jand g045(.dina(w_n117_1[2]),.dinb(w_n102_1[1]),.dout(n118),.clk(gclk));
	jnot g046(.din(Gic4),.dout(n119),.clk(gclk));
	jcb g047(.dina(w_n74_2[1]),.dinb(n119),.dout(n120));
	jxor g048(.dina(w_dff_B_nYQA3b499_0),.dinb(w_n93_0[0]),.dout(n121),.clk(gclk));
	jxor g049(.dina(w_Gid20_0[1]),.dinb(w_Gid16_0[1]),.dout(n122),.clk(gclk));
	jxor g050(.dina(w_Gid28_0[2]),.dinb(w_Gid24_0[2]),.dout(n123),.clk(gclk));
	jxor g051(.dina(n123),.dinb(n122),.dout(n124),.clk(gclk));
	jxor g052(.dina(n124),.dinb(w_n107_0[0]),.dout(n125),.clk(gclk));
	jxor g053(.dina(n125),.dinb(n121),.dout(n126),.clk(gclk));
	jnot g054(.din(w_n126_1[1]),.dout(n127),.clk(gclk));
	jnot g055(.din(Gic5),.dout(n128),.clk(gclk));
	jcb g056(.dina(w_n74_2[0]),.dinb(n128),.dout(n129));
	jxor g057(.dina(w_dff_B_ubnJPw2i5_0),.dinb(w_n97_0[0]),.dout(n130),.clk(gclk));
	jxor g058(.dina(w_Gid21_0[1]),.dinb(w_Gid17_0[1]),.dout(n131),.clk(gclk));
	jxor g059(.dina(w_Gid29_0[2]),.dinb(w_Gid25_0[2]),.dout(n132),.clk(gclk));
	jxor g060(.dina(n132),.dinb(n131),.dout(n133),.clk(gclk));
	jxor g061(.dina(n133),.dinb(w_n111_0[0]),.dout(n134),.clk(gclk));
	jxor g062(.dina(n134),.dinb(n130),.dout(n135),.clk(gclk));
	jand g063(.dina(w_n135_1[1]),.dinb(w_n127_1[2]),.dout(n136),.clk(gclk));
	jnot g064(.din(Gic1),.dout(n137),.clk(gclk));
	jcb g065(.dina(w_n74_1[2]),.dinb(n137),.dout(n138));
	jxor g066(.dina(w_Gid29_0[1]),.dinb(w_Gid28_0[1]),.dout(n139),.clk(gclk));
	jxor g067(.dina(w_Gid31_0[1]),.dinb(w_Gid30_0[1]),.dout(n140),.clk(gclk));
	jxor g068(.dina(n140),.dinb(n139),.dout(n141),.clk(gclk));
	jxor g069(.dina(w_n141_0[1]),.dinb(w_dff_B_fq2pqfIy1_1),.dout(n142),.clk(gclk));
	jxor g070(.dina(w_Gid25_0[1]),.dinb(w_Gid24_0[1]),.dout(n143),.clk(gclk));
	jxor g071(.dina(w_Gid27_0[1]),.dinb(w_Gid26_0[1]),.dout(n144),.clk(gclk));
	jxor g072(.dina(n144),.dinb(n143),.dout(n145),.clk(gclk));
	jxor g073(.dina(w_Gid5_0[1]),.dinb(w_Gid1_0[1]),.dout(n146),.clk(gclk));
	jxor g074(.dina(w_Gid13_0[1]),.dinb(w_Gid9_0[1]),.dout(n147),.clk(gclk));
	jxor g075(.dina(n147),.dinb(n146),.dout(n148),.clk(gclk));
	jxor g076(.dina(n148),.dinb(w_n145_0[1]),.dout(n149),.clk(gclk));
	jxor g077(.dina(n149),.dinb(n142),.dout(n150),.clk(gclk));
	jxor g078(.dina(w_n150_1[1]),.dinb(w_n87_1[0]),.dout(n151),.clk(gclk));
	jnot g079(.din(Gic3),.dout(n152),.clk(gclk));
	jcb g080(.dina(w_n74_1[1]),.dinb(n152),.dout(n153));
	jxor g081(.dina(w_dff_B_nOPe9sMB7_0),.dinb(w_n85_0[0]),.dout(n154),.clk(gclk));
	jxor g082(.dina(w_Gid7_0[1]),.dinb(w_Gid3_0[1]),.dout(n155),.clk(gclk));
	jxor g083(.dina(w_Gid15_0[1]),.dinb(w_Gid11_0[1]),.dout(n156),.clk(gclk));
	jxor g084(.dina(n156),.dinb(n155),.dout(n157),.clk(gclk));
	jxor g085(.dina(n157),.dinb(w_n141_0[0]),.dout(n158),.clk(gclk));
	jxor g086(.dina(n158),.dinb(n154),.dout(n159),.clk(gclk));
	jnot g087(.din(Gic2),.dout(n160),.clk(gclk));
	jcb g088(.dina(w_n74_1[0]),.dinb(n160),.dout(n161));
	jxor g089(.dina(w_dff_B_i2Mv9mSE2_0),.dinb(w_n78_0[0]),.dout(n162),.clk(gclk));
	jxor g090(.dina(w_Gid6_0[1]),.dinb(w_Gid2_0[1]),.dout(n163),.clk(gclk));
	jxor g091(.dina(w_Gid14_0[1]),.dinb(w_Gid10_0[1]),.dout(n164),.clk(gclk));
	jxor g092(.dina(n164),.dinb(n163),.dout(n165),.clk(gclk));
	jxor g093(.dina(n165),.dinb(w_n145_0[0]),.dout(n166),.clk(gclk));
	jxor g094(.dina(n166),.dinb(n162),.dout(n167),.clk(gclk));
	jand g095(.dina(w_n167_1[1]),.dinb(w_n159_1[1]),.dout(n168),.clk(gclk));
	jand g096(.dina(n168),.dinb(n151),.dout(n169),.clk(gclk));
	jxor g097(.dina(w_n167_1[0]),.dinb(w_n159_1[0]),.dout(n170),.clk(gclk));
	jand g098(.dina(w_n150_1[0]),.dinb(w_n87_0[2]),.dout(n171),.clk(gclk));
	jand g099(.dina(n171),.dinb(n170),.dout(n172),.clk(gclk));
	jcb g100(.dina(n172),.dinb(n169),.dout(n173));
	jand g101(.dina(w_n173_0[2]),.dinb(n136),.dout(n174),.clk(gclk));
	jand g102(.dina(w_n174_0[1]),.dinb(w_n118_0[1]),.dout(n175),.clk(gclk));
	jand g103(.dina(w_n175_1[1]),.dinb(w_n88_1[2]),.dout(n176),.clk(gclk));
	jxor g104(.dina(n176),.dinb(w_Gid0_0[0]),.dout(God0),.clk(gclk));
	jnot g105(.din(w_n150_0[2]),.dout(n178),.clk(gclk));
	jand g106(.dina(w_n175_1[0]),.dinb(w_n178_1[2]),.dout(n179),.clk(gclk));
	jxor g107(.dina(n179),.dinb(w_Gid1_0[0]),.dout(God1),.clk(gclk));
	jnot g108(.din(w_n167_0[2]),.dout(n181),.clk(gclk));
	jand g109(.dina(w_n175_0[2]),.dinb(w_n181_1[2]),.dout(n182),.clk(gclk));
	jxor g110(.dina(n182),.dinb(w_Gid2_0[0]),.dout(God2),.clk(gclk));
	jnot g111(.din(w_n159_0[2]),.dout(n184),.clk(gclk));
	jand g112(.dina(w_n175_0[1]),.dinb(w_n184_1[2]),.dout(n185),.clk(gclk));
	jxor g113(.dina(n185),.dinb(w_Gid3_0[0]),.dout(God3),.clk(gclk));
	jnot g114(.din(w_n102_1[0]),.dout(n187),.clk(gclk));
	jand g115(.dina(w_n116_1[0]),.dinb(w_n187_1[2]),.dout(n188),.clk(gclk));
	jand g116(.dina(w_n188_0[1]),.dinb(w_n174_0[0]),.dout(n189),.clk(gclk));
	jand g117(.dina(w_n189_1[1]),.dinb(w_n88_1[1]),.dout(n190),.clk(gclk));
	jxor g118(.dina(n190),.dinb(w_Gid4_0[0]),.dout(God4),.clk(gclk));
	jand g119(.dina(w_n189_1[0]),.dinb(w_n178_1[1]),.dout(n192),.clk(gclk));
	jxor g120(.dina(n192),.dinb(w_Gid5_0[0]),.dout(God5),.clk(gclk));
	jand g121(.dina(w_n189_0[2]),.dinb(w_n181_1[1]),.dout(n194),.clk(gclk));
	jxor g122(.dina(n194),.dinb(w_Gid6_0[0]),.dout(God6),.clk(gclk));
	jand g123(.dina(w_n189_0[1]),.dinb(w_n184_1[1]),.dout(n196),.clk(gclk));
	jxor g124(.dina(n196),.dinb(w_Gid7_0[0]),.dout(God7),.clk(gclk));
	jnot g125(.din(w_n135_1[0]),.dout(n198),.clk(gclk));
	jand g126(.dina(w_n198_1[2]),.dinb(w_n126_1[0]),.dout(n199),.clk(gclk));
	jand g127(.dina(w_n199_0[1]),.dinb(w_n118_0[0]),.dout(n200),.clk(gclk));
	jand g128(.dina(n200),.dinb(w_n173_0[1]),.dout(n201),.clk(gclk));
	jand g129(.dina(w_n201_1[1]),.dinb(w_n88_1[0]),.dout(n202),.clk(gclk));
	jxor g130(.dina(n202),.dinb(w_Gid8_0[0]),.dout(God8),.clk(gclk));
	jand g131(.dina(w_n201_1[0]),.dinb(w_n178_1[0]),.dout(n204),.clk(gclk));
	jxor g132(.dina(n204),.dinb(w_Gid9_0[0]),.dout(God9),.clk(gclk));
	jand g133(.dina(w_n201_0[2]),.dinb(w_n181_1[0]),.dout(n206),.clk(gclk));
	jxor g134(.dina(n206),.dinb(w_Gid10_0[0]),.dout(God10),.clk(gclk));
	jand g135(.dina(w_n201_0[1]),.dinb(w_n184_1[0]),.dout(n208),.clk(gclk));
	jxor g136(.dina(n208),.dinb(w_Gid11_0[0]),.dout(God11),.clk(gclk));
	jand g137(.dina(w_n199_0[0]),.dinb(w_n188_0[0]),.dout(n210),.clk(gclk));
	jand g138(.dina(n210),.dinb(w_n173_0[0]),.dout(n211),.clk(gclk));
	jand g139(.dina(w_n211_1[1]),.dinb(w_n88_0[2]),.dout(n212),.clk(gclk));
	jxor g140(.dina(n212),.dinb(w_Gid12_0[0]),.dout(God12),.clk(gclk));
	jand g141(.dina(w_n211_1[0]),.dinb(w_n178_0[2]),.dout(n214),.clk(gclk));
	jxor g142(.dina(n214),.dinb(w_Gid13_0[0]),.dout(God13),.clk(gclk));
	jand g143(.dina(w_n211_0[2]),.dinb(w_n181_0[2]),.dout(n216),.clk(gclk));
	jxor g144(.dina(n216),.dinb(w_Gid14_0[0]),.dout(God14),.clk(gclk));
	jand g145(.dina(w_n211_0[1]),.dinb(w_n184_0[2]),.dout(n218),.clk(gclk));
	jxor g146(.dina(n218),.dinb(w_Gid15_0[0]),.dout(God15),.clk(gclk));
	jand g147(.dina(w_n150_0[1]),.dinb(w_n88_0[1]),.dout(n220),.clk(gclk));
	jand g148(.dina(w_n181_0[1]),.dinb(w_n159_0[1]),.dout(n221),.clk(gclk));
	jxor g149(.dina(w_n116_0[2]),.dinb(w_n102_0[2]),.dout(n222),.clk(gclk));
	jand g150(.dina(w_n135_0[2]),.dinb(w_n126_0[2]),.dout(n223),.clk(gclk));
	jand g151(.dina(n223),.dinb(n222),.dout(n224),.clk(gclk));
	jxor g152(.dina(w_n135_0[1]),.dinb(w_n126_0[1]),.dout(n225),.clk(gclk));
	jand g153(.dina(w_n116_0[1]),.dinb(w_n102_0[1]),.dout(n226),.clk(gclk));
	jand g154(.dina(n226),.dinb(n225),.dout(n227),.clk(gclk));
	jcb g155(.dina(n227),.dinb(n224),.dout(n228));
	jand g156(.dina(w_n228_0[1]),.dinb(n221),.dout(n229),.clk(gclk));
	jand g157(.dina(w_n229_0[1]),.dinb(w_n220_0[1]),.dout(n230),.clk(gclk));
	jand g158(.dina(w_n230_1[1]),.dinb(w_n127_1[1]),.dout(n231),.clk(gclk));
	jxor g159(.dina(n231),.dinb(w_Gid16_0[0]),.dout(God16),.clk(gclk));
	jand g160(.dina(w_n230_1[0]),.dinb(w_n198_1[1]),.dout(n233),.clk(gclk));
	jxor g161(.dina(n233),.dinb(w_Gid17_0[0]),.dout(God17),.clk(gclk));
	jand g162(.dina(w_n230_0[2]),.dinb(w_n117_1[1]),.dout(n235),.clk(gclk));
	jxor g163(.dina(n235),.dinb(w_Gid18_0[0]),.dout(God18),.clk(gclk));
	jand g164(.dina(w_n230_0[1]),.dinb(w_n187_1[1]),.dout(n237),.clk(gclk));
	jxor g165(.dina(n237),.dinb(w_Gid19_0[0]),.dout(God19),.clk(gclk));
	jand g166(.dina(w_n167_0[1]),.dinb(w_n184_0[1]),.dout(n239),.clk(gclk));
	jand g167(.dina(w_n228_0[0]),.dinb(n239),.dout(n240),.clk(gclk));
	jand g168(.dina(w_n240_0[1]),.dinb(w_n220_0[0]),.dout(n241),.clk(gclk));
	jand g169(.dina(w_n241_1[1]),.dinb(w_n127_1[0]),.dout(n242),.clk(gclk));
	jxor g170(.dina(n242),.dinb(w_Gid20_0[0]),.dout(God20),.clk(gclk));
	jand g171(.dina(w_n241_1[0]),.dinb(w_n198_1[0]),.dout(n244),.clk(gclk));
	jxor g172(.dina(n244),.dinb(w_Gid21_0[0]),.dout(God21),.clk(gclk));
	jand g173(.dina(w_n241_0[2]),.dinb(w_n117_1[0]),.dout(n246),.clk(gclk));
	jxor g174(.dina(n246),.dinb(w_Gid22_0[0]),.dout(God22),.clk(gclk));
	jand g175(.dina(w_n241_0[1]),.dinb(w_n187_1[0]),.dout(n248),.clk(gclk));
	jxor g176(.dina(n248),.dinb(w_Gid23_0[0]),.dout(God23),.clk(gclk));
	jand g177(.dina(w_n178_0[1]),.dinb(w_n87_0[1]),.dout(n250),.clk(gclk));
	jand g178(.dina(w_n229_0[0]),.dinb(w_n250_0[1]),.dout(n251),.clk(gclk));
	jand g179(.dina(w_n251_1[1]),.dinb(w_n127_0[2]),.dout(n252),.clk(gclk));
	jxor g180(.dina(n252),.dinb(w_Gid24_0[0]),.dout(God24),.clk(gclk));
	jand g181(.dina(w_n251_1[0]),.dinb(w_n198_0[2]),.dout(n254),.clk(gclk));
	jxor g182(.dina(n254),.dinb(w_Gid25_0[0]),.dout(God25),.clk(gclk));
	jand g183(.dina(w_n251_0[2]),.dinb(w_n117_0[2]),.dout(n256),.clk(gclk));
	jxor g184(.dina(n256),.dinb(w_Gid26_0[0]),.dout(God26),.clk(gclk));
	jand g185(.dina(w_n251_0[1]),.dinb(w_n187_0[2]),.dout(n258),.clk(gclk));
	jxor g186(.dina(n258),.dinb(w_Gid27_0[0]),.dout(God27),.clk(gclk));
	jand g187(.dina(w_n240_0[0]),.dinb(w_n250_0[0]),.dout(n260),.clk(gclk));
	jand g188(.dina(w_n260_1[1]),.dinb(w_n127_0[1]),.dout(n261),.clk(gclk));
	jxor g189(.dina(n261),.dinb(w_Gid28_0[0]),.dout(God28),.clk(gclk));
	jand g190(.dina(w_n260_1[0]),.dinb(w_n198_0[1]),.dout(n263),.clk(gclk));
	jxor g191(.dina(n263),.dinb(w_Gid29_0[0]),.dout(God29),.clk(gclk));
	jand g192(.dina(w_n260_0[2]),.dinb(w_n117_0[1]),.dout(n265),.clk(gclk));
	jxor g193(.dina(n265),.dinb(w_Gid30_0[0]),.dout(God30),.clk(gclk));
	jand g194(.dina(w_n260_0[1]),.dinb(w_n187_0[1]),.dout(n267),.clk(gclk));
	jxor g195(.dina(n267),.dinb(w_Gid31_0[0]),.dout(God31),.clk(gclk));
	jspl3 jspl3_w_Gid0_0(.douta(w_dff_A_jeIqdny36_0),.doutb(w_Gid0_0[1]),.doutc(w_Gid0_0[2]),.din(Gid0));
	jspl3 jspl3_w_Gid1_0(.douta(w_dff_A_ibDwxNCx3_0),.doutb(w_Gid1_0[1]),.doutc(w_Gid1_0[2]),.din(Gid1));
	jspl3 jspl3_w_Gid2_0(.douta(w_dff_A_asTtwopN9_0),.doutb(w_Gid2_0[1]),.doutc(w_Gid2_0[2]),.din(Gid2));
	jspl3 jspl3_w_Gid3_0(.douta(w_dff_A_jJuM7kdD5_0),.doutb(w_Gid3_0[1]),.doutc(w_Gid3_0[2]),.din(Gid3));
	jspl3 jspl3_w_Gid4_0(.douta(w_dff_A_D8w0sMRT0_0),.doutb(w_Gid4_0[1]),.doutc(w_Gid4_0[2]),.din(Gid4));
	jspl3 jspl3_w_Gid5_0(.douta(w_dff_A_f4JIbIaN0_0),.doutb(w_Gid5_0[1]),.doutc(w_Gid5_0[2]),.din(Gid5));
	jspl3 jspl3_w_Gid6_0(.douta(w_dff_A_7fxMyzXe9_0),.doutb(w_Gid6_0[1]),.doutc(w_Gid6_0[2]),.din(Gid6));
	jspl3 jspl3_w_Gid7_0(.douta(w_dff_A_DMwycXsd8_0),.doutb(w_Gid7_0[1]),.doutc(w_Gid7_0[2]),.din(Gid7));
	jspl3 jspl3_w_Gid8_0(.douta(w_dff_A_Fm81bVXb4_0),.doutb(w_Gid8_0[1]),.doutc(w_Gid8_0[2]),.din(Gid8));
	jspl3 jspl3_w_Gid9_0(.douta(w_dff_A_KnxHH5LI4_0),.doutb(w_Gid9_0[1]),.doutc(w_Gid9_0[2]),.din(Gid9));
	jspl3 jspl3_w_Gid10_0(.douta(w_dff_A_J2bJJcFI8_0),.doutb(w_Gid10_0[1]),.doutc(w_Gid10_0[2]),.din(Gid10));
	jspl3 jspl3_w_Gid11_0(.douta(w_dff_A_Lni5NrPW5_0),.doutb(w_Gid11_0[1]),.doutc(w_Gid11_0[2]),.din(Gid11));
	jspl3 jspl3_w_Gid12_0(.douta(w_dff_A_1YGnxI0q7_0),.doutb(w_Gid12_0[1]),.doutc(w_Gid12_0[2]),.din(Gid12));
	jspl3 jspl3_w_Gid13_0(.douta(w_dff_A_iv4e9N5q4_0),.doutb(w_Gid13_0[1]),.doutc(w_Gid13_0[2]),.din(Gid13));
	jspl3 jspl3_w_Gid14_0(.douta(w_dff_A_QIjOxqaN9_0),.doutb(w_Gid14_0[1]),.doutc(w_Gid14_0[2]),.din(Gid14));
	jspl3 jspl3_w_Gid15_0(.douta(w_dff_A_4KrvNnKl3_0),.doutb(w_Gid15_0[1]),.doutc(w_Gid15_0[2]),.din(Gid15));
	jspl3 jspl3_w_Gid16_0(.douta(w_dff_A_7a90pXgD9_0),.doutb(w_Gid16_0[1]),.doutc(w_Gid16_0[2]),.din(Gid16));
	jspl3 jspl3_w_Gid17_0(.douta(w_dff_A_TLDVzjjS5_0),.doutb(w_Gid17_0[1]),.doutc(w_Gid17_0[2]),.din(Gid17));
	jspl3 jspl3_w_Gid18_0(.douta(w_dff_A_pEGxduJo7_0),.doutb(w_Gid18_0[1]),.doutc(w_Gid18_0[2]),.din(Gid18));
	jspl3 jspl3_w_Gid19_0(.douta(w_dff_A_nCnJAGQY6_0),.doutb(w_Gid19_0[1]),.doutc(w_Gid19_0[2]),.din(Gid19));
	jspl3 jspl3_w_Gid20_0(.douta(w_dff_A_8AF4rwWG4_0),.doutb(w_Gid20_0[1]),.doutc(w_Gid20_0[2]),.din(Gid20));
	jspl3 jspl3_w_Gid21_0(.douta(w_dff_A_SBxBORC27_0),.doutb(w_Gid21_0[1]),.doutc(w_Gid21_0[2]),.din(Gid21));
	jspl3 jspl3_w_Gid22_0(.douta(w_dff_A_ZlF6DRNS8_0),.doutb(w_Gid22_0[1]),.doutc(w_Gid22_0[2]),.din(Gid22));
	jspl3 jspl3_w_Gid23_0(.douta(w_dff_A_PiQJmDTh0_0),.doutb(w_Gid23_0[1]),.doutc(w_Gid23_0[2]),.din(Gid23));
	jspl3 jspl3_w_Gid24_0(.douta(w_dff_A_2bZYM1jj9_0),.doutb(w_Gid24_0[1]),.doutc(w_Gid24_0[2]),.din(Gid24));
	jspl3 jspl3_w_Gid25_0(.douta(w_dff_A_p0JsYRz87_0),.doutb(w_Gid25_0[1]),.doutc(w_Gid25_0[2]),.din(Gid25));
	jspl3 jspl3_w_Gid26_0(.douta(w_dff_A_mLEMYJRM9_0),.doutb(w_Gid26_0[1]),.doutc(w_Gid26_0[2]),.din(Gid26));
	jspl3 jspl3_w_Gid27_0(.douta(w_dff_A_atPkpVhr5_0),.doutb(w_Gid27_0[1]),.doutc(w_Gid27_0[2]),.din(Gid27));
	jspl3 jspl3_w_Gid28_0(.douta(w_dff_A_KqvraJus8_0),.doutb(w_Gid28_0[1]),.doutc(w_Gid28_0[2]),.din(Gid28));
	jspl3 jspl3_w_Gid29_0(.douta(w_dff_A_lpdSTX472_0),.doutb(w_Gid29_0[1]),.doutc(w_Gid29_0[2]),.din(Gid29));
	jspl3 jspl3_w_Gid30_0(.douta(w_dff_A_PGuNR5kM5_0),.doutb(w_Gid30_0[1]),.doutc(w_Gid30_0[2]),.din(Gid30));
	jspl3 jspl3_w_Gid31_0(.douta(w_dff_A_Mk7fOtus9_0),.doutb(w_Gid31_0[1]),.doutc(w_Gid31_0[2]),.din(Gid31));
	jspl3 jspl3_w_n74_0(.douta(w_n74_0[0]),.doutb(w_n74_0[1]),.doutc(w_n74_0[2]),.din(n74));
	jspl3 jspl3_w_n74_1(.douta(w_n74_1[0]),.doutb(w_n74_1[1]),.doutc(w_n74_1[2]),.din(w_n74_0[0]));
	jspl3 jspl3_w_n74_2(.douta(w_n74_2[0]),.doutb(w_n74_2[1]),.doutc(w_n74_2[2]),.din(w_n74_0[1]));
	jspl jspl_w_n74_3(.douta(w_n74_3[0]),.doutb(w_n74_3[1]),.din(w_n74_0[2]));
	jspl jspl_w_n78_0(.douta(w_n78_0[0]),.doutb(w_n78_0[1]),.din(n78));
	jspl jspl_w_n85_0(.douta(w_n85_0[0]),.doutb(w_n85_0[1]),.din(n85));
	jspl3 jspl3_w_n87_0(.douta(w_n87_0[0]),.doutb(w_dff_A_PXTVRGeM9_1),.doutc(w_n87_0[2]),.din(n87));
	jspl jspl_w_n87_1(.douta(w_n87_1[0]),.doutb(w_n87_1[1]),.din(w_n87_0[0]));
	jspl3 jspl3_w_n88_0(.douta(w_dff_A_7HOZnrRL8_0),.doutb(w_n88_0[1]),.doutc(w_dff_A_cMWeQ5XI8_2),.din(n88));
	jspl3 jspl3_w_n88_1(.douta(w_n88_1[0]),.doutb(w_n88_1[1]),.doutc(w_n88_1[2]),.din(w_n88_0[0]));
	jspl jspl_w_n93_0(.douta(w_n93_0[0]),.doutb(w_n93_0[1]),.din(n93));
	jspl jspl_w_n97_0(.douta(w_n97_0[0]),.doutb(w_n97_0[1]),.din(n97));
	jspl3 jspl3_w_n102_0(.douta(w_n102_0[0]),.doutb(w_n102_0[1]),.doutc(w_n102_0[2]),.din(n102));
	jspl jspl_w_n102_1(.douta(w_n102_1[0]),.doutb(w_dff_A_onFBGz5h5_1),.din(w_n102_0[0]));
	jspl jspl_w_n107_0(.douta(w_n107_0[0]),.doutb(w_n107_0[1]),.din(n107));
	jspl jspl_w_n111_0(.douta(w_n111_0[0]),.doutb(w_n111_0[1]),.din(n111));
	jspl3 jspl3_w_n116_0(.douta(w_n116_0[0]),.doutb(w_n116_0[1]),.doutc(w_n116_0[2]),.din(n116));
	jspl jspl_w_n116_1(.douta(w_dff_A_QG81S6Au8_0),.doutb(w_n116_1[1]),.din(w_n116_0[0]));
	jspl3 jspl3_w_n117_0(.douta(w_n117_0[0]),.doutb(w_dff_A_VJiCPsNs4_1),.doutc(w_dff_A_umK8VC3f9_2),.din(n117));
	jspl3 jspl3_w_n117_1(.douta(w_dff_A_RdyzR5Yi3_0),.doutb(w_dff_A_k5aMHF8R6_1),.doutc(w_n117_1[2]),.din(w_n117_0[0]));
	jspl jspl_w_n118_0(.douta(w_n118_0[0]),.doutb(w_dff_A_Gay8MZ4x5_1),.din(n118));
	jspl3 jspl3_w_n126_0(.douta(w_n126_0[0]),.doutb(w_n126_0[1]),.doutc(w_n126_0[2]),.din(n126));
	jspl jspl_w_n126_1(.douta(w_dff_A_6fvZ8SAh2_0),.doutb(w_n126_1[1]),.din(w_n126_0[0]));
	jspl3 jspl3_w_n127_0(.douta(w_n127_0[0]),.doutb(w_dff_A_QP3bYQP69_1),.doutc(w_dff_A_jozhULJA9_2),.din(n127));
	jspl3 jspl3_w_n127_1(.douta(w_dff_A_iUsVz9Of4_0),.doutb(w_dff_A_AFC26J8h4_1),.doutc(w_n127_1[2]),.din(w_n127_0[0]));
	jspl3 jspl3_w_n135_0(.douta(w_n135_0[0]),.doutb(w_n135_0[1]),.doutc(w_n135_0[2]),.din(n135));
	jspl jspl_w_n135_1(.douta(w_n135_1[0]),.doutb(w_dff_A_o7MXsCVg9_1),.din(w_n135_0[0]));
	jspl jspl_w_n141_0(.douta(w_n141_0[0]),.doutb(w_n141_0[1]),.din(n141));
	jspl jspl_w_n145_0(.douta(w_n145_0[0]),.doutb(w_n145_0[1]),.din(n145));
	jspl3 jspl3_w_n150_0(.douta(w_n150_0[0]),.doutb(w_dff_A_7VTeUlZZ6_1),.doutc(w_n150_0[2]),.din(n150));
	jspl jspl_w_n150_1(.douta(w_n150_1[0]),.doutb(w_n150_1[1]),.din(w_n150_0[0]));
	jspl3 jspl3_w_n159_0(.douta(w_n159_0[0]),.doutb(w_dff_A_USYzVecP0_1),.doutc(w_n159_0[2]),.din(n159));
	jspl jspl_w_n159_1(.douta(w_n159_1[0]),.doutb(w_n159_1[1]),.din(w_n159_0[0]));
	jspl3 jspl3_w_n167_0(.douta(w_n167_0[0]),.doutb(w_dff_A_ZwEhqkxI7_1),.doutc(w_n167_0[2]),.din(n167));
	jspl jspl_w_n167_1(.douta(w_n167_1[0]),.doutb(w_n167_1[1]),.din(w_n167_0[0]));
	jspl3 jspl3_w_n173_0(.douta(w_dff_A_nkkr6ssB2_0),.doutb(w_dff_A_SoPSj0JI0_1),.doutc(w_n173_0[2]),.din(n173));
	jspl jspl_w_n174_0(.douta(w_n174_0[0]),.doutb(w_n174_0[1]),.din(n174));
	jspl3 jspl3_w_n175_0(.douta(w_n175_0[0]),.doutb(w_n175_0[1]),.doutc(w_n175_0[2]),.din(n175));
	jspl jspl_w_n175_1(.douta(w_n175_1[0]),.doutb(w_n175_1[1]),.din(w_n175_0[0]));
	jspl3 jspl3_w_n178_0(.douta(w_dff_A_d3Pa53nW2_0),.doutb(w_n178_0[1]),.doutc(w_dff_A_vdMCMSdo5_2),.din(n178));
	jspl3 jspl3_w_n178_1(.douta(w_n178_1[0]),.doutb(w_n178_1[1]),.doutc(w_n178_1[2]),.din(w_n178_0[0]));
	jspl3 jspl3_w_n181_0(.douta(w_dff_A_TSdGAzNV8_0),.doutb(w_n181_0[1]),.doutc(w_dff_A_JArBfUQ79_2),.din(n181));
	jspl3 jspl3_w_n181_1(.douta(w_n181_1[0]),.doutb(w_n181_1[1]),.doutc(w_n181_1[2]),.din(w_n181_0[0]));
	jspl3 jspl3_w_n184_0(.douta(w_dff_A_WhzBcMHk9_0),.doutb(w_n184_0[1]),.doutc(w_dff_A_F0a4qMEL1_2),.din(n184));
	jspl3 jspl3_w_n184_1(.douta(w_n184_1[0]),.doutb(w_n184_1[1]),.doutc(w_n184_1[2]),.din(w_n184_0[0]));
	jspl3 jspl3_w_n187_0(.douta(w_n187_0[0]),.doutb(w_dff_A_5g65sS2q0_1),.doutc(w_dff_A_SI7LRVvI5_2),.din(n187));
	jspl3 jspl3_w_n187_1(.douta(w_dff_A_WAcsnX4T5_0),.doutb(w_dff_A_cru1nvzF8_1),.doutc(w_n187_1[2]),.din(w_n187_0[0]));
	jspl jspl_w_n188_0(.douta(w_n188_0[0]),.doutb(w_dff_A_8UoaUcmQ7_1),.din(n188));
	jspl3 jspl3_w_n189_0(.douta(w_n189_0[0]),.doutb(w_n189_0[1]),.doutc(w_n189_0[2]),.din(n189));
	jspl jspl_w_n189_1(.douta(w_n189_1[0]),.doutb(w_n189_1[1]),.din(w_n189_0[0]));
	jspl3 jspl3_w_n198_0(.douta(w_n198_0[0]),.doutb(w_dff_A_wxGtXfff4_1),.doutc(w_dff_A_I8uXnHgx3_2),.din(n198));
	jspl3 jspl3_w_n198_1(.douta(w_dff_A_obfMM42W9_0),.doutb(w_dff_A_ybqClvk39_1),.doutc(w_n198_1[2]),.din(w_n198_0[0]));
	jspl jspl_w_n199_0(.douta(w_n199_0[0]),.doutb(w_n199_0[1]),.din(n199));
	jspl3 jspl3_w_n201_0(.douta(w_n201_0[0]),.doutb(w_n201_0[1]),.doutc(w_n201_0[2]),.din(n201));
	jspl jspl_w_n201_1(.douta(w_n201_1[0]),.doutb(w_n201_1[1]),.din(w_n201_0[0]));
	jspl3 jspl3_w_n211_0(.douta(w_n211_0[0]),.doutb(w_n211_0[1]),.doutc(w_n211_0[2]),.din(n211));
	jspl jspl_w_n211_1(.douta(w_n211_1[0]),.doutb(w_n211_1[1]),.din(w_n211_0[0]));
	jspl jspl_w_n220_0(.douta(w_n220_0[0]),.doutb(w_n220_0[1]),.din(w_dff_B_ZNirXdbH6_2));
	jspl jspl_w_n228_0(.douta(w_n228_0[0]),.doutb(w_n228_0[1]),.din(n228));
	jspl jspl_w_n229_0(.douta(w_n229_0[0]),.doutb(w_n229_0[1]),.din(n229));
	jspl3 jspl3_w_n230_0(.douta(w_n230_0[0]),.doutb(w_n230_0[1]),.doutc(w_n230_0[2]),.din(n230));
	jspl jspl_w_n230_1(.douta(w_n230_1[0]),.doutb(w_n230_1[1]),.din(w_n230_0[0]));
	jspl jspl_w_n240_0(.douta(w_n240_0[0]),.doutb(w_n240_0[1]),.din(n240));
	jspl3 jspl3_w_n241_0(.douta(w_n241_0[0]),.doutb(w_n241_0[1]),.doutc(w_n241_0[2]),.din(n241));
	jspl jspl_w_n241_1(.douta(w_n241_1[0]),.doutb(w_n241_1[1]),.din(w_n241_0[0]));
	jspl jspl_w_n250_0(.douta(w_n250_0[0]),.doutb(w_n250_0[1]),.din(w_dff_B_UC88yyfr6_2));
	jspl3 jspl3_w_n251_0(.douta(w_n251_0[0]),.doutb(w_n251_0[1]),.doutc(w_n251_0[2]),.din(n251));
	jspl jspl_w_n251_1(.douta(w_n251_1[0]),.doutb(w_n251_1[1]),.din(w_n251_0[0]));
	jspl3 jspl3_w_n260_0(.douta(w_n260_0[0]),.doutb(w_n260_0[1]),.doutc(w_n260_0[2]),.din(n260));
	jspl jspl_w_n260_1(.douta(w_n260_1[0]),.doutb(w_n260_1[1]),.din(w_n260_0[0]));
	jdff dff_A_Gay8MZ4x5_1(.dout(w_n118_0[1]),.din(w_dff_A_Gay8MZ4x5_1),.clk(gclk));
	jdff dff_A_8UoaUcmQ7_1(.dout(w_n188_0[1]),.din(w_dff_A_8UoaUcmQ7_1),.clk(gclk));
	jdff dff_A_nkkr6ssB2_0(.dout(w_n173_0[0]),.din(w_dff_A_nkkr6ssB2_0),.clk(gclk));
	jdff dff_A_SoPSj0JI0_1(.dout(w_n173_0[1]),.din(w_dff_A_SoPSj0JI0_1),.clk(gclk));
	jdff dff_A_z8wTnRGS4_0(.dout(w_n127_1[0]),.din(w_dff_A_z8wTnRGS4_0),.clk(gclk));
	jdff dff_A_p0OCm6EC3_0(.dout(w_dff_A_z8wTnRGS4_0),.din(w_dff_A_p0OCm6EC3_0),.clk(gclk));
	jdff dff_A_iUsVz9Of4_0(.dout(w_dff_A_p0OCm6EC3_0),.din(w_dff_A_iUsVz9Of4_0),.clk(gclk));
	jdff dff_A_D2t15BiB9_1(.dout(w_n127_1[1]),.din(w_dff_A_D2t15BiB9_1),.clk(gclk));
	jdff dff_A_VvqVNZHs2_1(.dout(w_dff_A_D2t15BiB9_1),.din(w_dff_A_VvqVNZHs2_1),.clk(gclk));
	jdff dff_A_AFC26J8h4_1(.dout(w_dff_A_VvqVNZHs2_1),.din(w_dff_A_AFC26J8h4_1),.clk(gclk));
	jdff dff_A_gL4MMgIh2_0(.dout(w_n198_1[0]),.din(w_dff_A_gL4MMgIh2_0),.clk(gclk));
	jdff dff_A_VflmckS26_0(.dout(w_dff_A_gL4MMgIh2_0),.din(w_dff_A_VflmckS26_0),.clk(gclk));
	jdff dff_A_obfMM42W9_0(.dout(w_dff_A_VflmckS26_0),.din(w_dff_A_obfMM42W9_0),.clk(gclk));
	jdff dff_A_WxCg7RGe8_1(.dout(w_n198_1[1]),.din(w_dff_A_WxCg7RGe8_1),.clk(gclk));
	jdff dff_A_dVq2s78T0_1(.dout(w_dff_A_WxCg7RGe8_1),.din(w_dff_A_dVq2s78T0_1),.clk(gclk));
	jdff dff_A_ybqClvk39_1(.dout(w_dff_A_dVq2s78T0_1),.din(w_dff_A_ybqClvk39_1),.clk(gclk));
	jdff dff_A_mlZA7mzT3_0(.dout(w_n117_1[0]),.din(w_dff_A_mlZA7mzT3_0),.clk(gclk));
	jdff dff_A_m3AhxUKP9_0(.dout(w_dff_A_mlZA7mzT3_0),.din(w_dff_A_m3AhxUKP9_0),.clk(gclk));
	jdff dff_A_RdyzR5Yi3_0(.dout(w_dff_A_m3AhxUKP9_0),.din(w_dff_A_RdyzR5Yi3_0),.clk(gclk));
	jdff dff_A_lfU4Xgec4_1(.dout(w_n117_1[1]),.din(w_dff_A_lfU4Xgec4_1),.clk(gclk));
	jdff dff_A_E0PG8tGi1_1(.dout(w_dff_A_lfU4Xgec4_1),.din(w_dff_A_E0PG8tGi1_1),.clk(gclk));
	jdff dff_A_k5aMHF8R6_1(.dout(w_dff_A_E0PG8tGi1_1),.din(w_dff_A_k5aMHF8R6_1),.clk(gclk));
	jdff dff_B_ZNirXdbH6_2(.din(n220),.dout(w_dff_B_ZNirXdbH6_2),.clk(gclk));
	jdff dff_A_j4XMoKDy1_0(.dout(w_n88_0[0]),.din(w_dff_A_j4XMoKDy1_0),.clk(gclk));
	jdff dff_A_gfYr5qa00_0(.dout(w_dff_A_j4XMoKDy1_0),.din(w_dff_A_gfYr5qa00_0),.clk(gclk));
	jdff dff_A_7HOZnrRL8_0(.dout(w_dff_A_gfYr5qa00_0),.din(w_dff_A_7HOZnrRL8_0),.clk(gclk));
	jdff dff_A_a0CkAKZ58_2(.dout(w_n88_0[2]),.din(w_dff_A_a0CkAKZ58_2),.clk(gclk));
	jdff dff_A_we2xVxLm6_2(.dout(w_dff_A_a0CkAKZ58_2),.din(w_dff_A_we2xVxLm6_2),.clk(gclk));
	jdff dff_A_cMWeQ5XI8_2(.dout(w_dff_A_we2xVxLm6_2),.din(w_dff_A_cMWeQ5XI8_2),.clk(gclk));
	jdff dff_A_zKjvttGZ3_0(.dout(w_n187_1[0]),.din(w_dff_A_zKjvttGZ3_0),.clk(gclk));
	jdff dff_A_xNDejBvk0_0(.dout(w_dff_A_zKjvttGZ3_0),.din(w_dff_A_xNDejBvk0_0),.clk(gclk));
	jdff dff_A_WAcsnX4T5_0(.dout(w_dff_A_xNDejBvk0_0),.din(w_dff_A_WAcsnX4T5_0),.clk(gclk));
	jdff dff_A_MLKUktyu2_1(.dout(w_n187_1[1]),.din(w_dff_A_MLKUktyu2_1),.clk(gclk));
	jdff dff_A_mZ7wmJHc4_1(.dout(w_dff_A_MLKUktyu2_1),.din(w_dff_A_mZ7wmJHc4_1),.clk(gclk));
	jdff dff_A_cru1nvzF8_1(.dout(w_dff_A_mZ7wmJHc4_1),.din(w_dff_A_cru1nvzF8_1),.clk(gclk));
	jdff dff_A_t8diCatx3_0(.dout(w_n181_0[0]),.din(w_dff_A_t8diCatx3_0),.clk(gclk));
	jdff dff_A_FEisqJMX8_0(.dout(w_dff_A_t8diCatx3_0),.din(w_dff_A_FEisqJMX8_0),.clk(gclk));
	jdff dff_A_TSdGAzNV8_0(.dout(w_dff_A_FEisqJMX8_0),.din(w_dff_A_TSdGAzNV8_0),.clk(gclk));
	jdff dff_A_MAsuxIbO7_2(.dout(w_n181_0[2]),.din(w_dff_A_MAsuxIbO7_2),.clk(gclk));
	jdff dff_A_3T3QLBvE1_2(.dout(w_dff_A_MAsuxIbO7_2),.din(w_dff_A_3T3QLBvE1_2),.clk(gclk));
	jdff dff_A_JArBfUQ79_2(.dout(w_dff_A_3T3QLBvE1_2),.din(w_dff_A_JArBfUQ79_2),.clk(gclk));
	jdff dff_A_vio35cWh5_1(.dout(w_n127_0[1]),.din(w_dff_A_vio35cWh5_1),.clk(gclk));
	jdff dff_A_36jn2a659_1(.dout(w_dff_A_vio35cWh5_1),.din(w_dff_A_36jn2a659_1),.clk(gclk));
	jdff dff_A_QP3bYQP69_1(.dout(w_dff_A_36jn2a659_1),.din(w_dff_A_QP3bYQP69_1),.clk(gclk));
	jdff dff_A_g3WR95nz3_2(.dout(w_n127_0[2]),.din(w_dff_A_g3WR95nz3_2),.clk(gclk));
	jdff dff_A_jkOEhk0c1_2(.dout(w_dff_A_g3WR95nz3_2),.din(w_dff_A_jkOEhk0c1_2),.clk(gclk));
	jdff dff_A_jozhULJA9_2(.dout(w_dff_A_jkOEhk0c1_2),.din(w_dff_A_jozhULJA9_2),.clk(gclk));
	jdff dff_A_6fvZ8SAh2_0(.dout(w_n126_1[0]),.din(w_dff_A_6fvZ8SAh2_0),.clk(gclk));
	jdff dff_A_GQdN42S37_1(.dout(w_n198_0[1]),.din(w_dff_A_GQdN42S37_1),.clk(gclk));
	jdff dff_A_FOg1v7fp9_1(.dout(w_dff_A_GQdN42S37_1),.din(w_dff_A_FOg1v7fp9_1),.clk(gclk));
	jdff dff_A_wxGtXfff4_1(.dout(w_dff_A_FOg1v7fp9_1),.din(w_dff_A_wxGtXfff4_1),.clk(gclk));
	jdff dff_A_iJoDg3Ir3_2(.dout(w_n198_0[2]),.din(w_dff_A_iJoDg3Ir3_2),.clk(gclk));
	jdff dff_A_C72QquDl7_2(.dout(w_dff_A_iJoDg3Ir3_2),.din(w_dff_A_C72QquDl7_2),.clk(gclk));
	jdff dff_A_I8uXnHgx3_2(.dout(w_dff_A_C72QquDl7_2),.din(w_dff_A_I8uXnHgx3_2),.clk(gclk));
	jdff dff_A_o7MXsCVg9_1(.dout(w_n135_1[1]),.din(w_dff_A_o7MXsCVg9_1),.clk(gclk));
	jdff dff_A_ohslviSy4_1(.dout(w_n117_0[1]),.din(w_dff_A_ohslviSy4_1),.clk(gclk));
	jdff dff_A_uB2Dc9v70_1(.dout(w_dff_A_ohslviSy4_1),.din(w_dff_A_uB2Dc9v70_1),.clk(gclk));
	jdff dff_A_VJiCPsNs4_1(.dout(w_dff_A_uB2Dc9v70_1),.din(w_dff_A_VJiCPsNs4_1),.clk(gclk));
	jdff dff_A_ONG3ilCy9_2(.dout(w_n117_0[2]),.din(w_dff_A_ONG3ilCy9_2),.clk(gclk));
	jdff dff_A_bmfCiTBG4_2(.dout(w_dff_A_ONG3ilCy9_2),.din(w_dff_A_bmfCiTBG4_2),.clk(gclk));
	jdff dff_A_umK8VC3f9_2(.dout(w_dff_A_bmfCiTBG4_2),.din(w_dff_A_umK8VC3f9_2),.clk(gclk));
	jdff dff_A_QG81S6Au8_0(.dout(w_n116_1[0]),.din(w_dff_A_QG81S6Au8_0),.clk(gclk));
	jdff dff_B_ubnJPw2i5_0(.din(n129),.dout(w_dff_B_ubnJPw2i5_0),.clk(gclk));
	jdff dff_B_nYQA3b499_0(.din(n120),.dout(w_dff_B_nYQA3b499_0),.clk(gclk));
	jdff dff_B_qL0lohj90_1(.din(n104),.dout(w_dff_B_qL0lohj90_1),.clk(gclk));
	jdff dff_A_ZwEhqkxI7_1(.dout(w_n167_0[1]),.din(w_dff_A_ZwEhqkxI7_1),.clk(gclk));
	jdff dff_A_4NXxozkh3_0(.dout(w_Gid10_0[0]),.din(w_dff_A_4NXxozkh3_0),.clk(gclk));
	jdff dff_A_Lr87YYC90_0(.dout(w_dff_A_4NXxozkh3_0),.din(w_dff_A_Lr87YYC90_0),.clk(gclk));
	jdff dff_A_8yOhhC1f0_0(.dout(w_dff_A_Lr87YYC90_0),.din(w_dff_A_8yOhhC1f0_0),.clk(gclk));
	jdff dff_A_M1h9aFMj4_0(.dout(w_dff_A_8yOhhC1f0_0),.din(w_dff_A_M1h9aFMj4_0),.clk(gclk));
	jdff dff_A_i9j5lDzb9_0(.dout(w_dff_A_M1h9aFMj4_0),.din(w_dff_A_i9j5lDzb9_0),.clk(gclk));
	jdff dff_A_vGfJnd7g9_0(.dout(w_dff_A_i9j5lDzb9_0),.din(w_dff_A_vGfJnd7g9_0),.clk(gclk));
	jdff dff_A_do0Lp34X4_0(.dout(w_dff_A_vGfJnd7g9_0),.din(w_dff_A_do0Lp34X4_0),.clk(gclk));
	jdff dff_A_bqk6m5BF1_0(.dout(w_dff_A_do0Lp34X4_0),.din(w_dff_A_bqk6m5BF1_0),.clk(gclk));
	jdff dff_A_J2bJJcFI8_0(.dout(w_dff_A_bqk6m5BF1_0),.din(w_dff_A_J2bJJcFI8_0),.clk(gclk));
	jdff dff_A_Y7lcpacD6_0(.dout(w_Gid2_0[0]),.din(w_dff_A_Y7lcpacD6_0),.clk(gclk));
	jdff dff_A_hhVzoZaR9_0(.dout(w_dff_A_Y7lcpacD6_0),.din(w_dff_A_hhVzoZaR9_0),.clk(gclk));
	jdff dff_A_P6cRG2mZ2_0(.dout(w_dff_A_hhVzoZaR9_0),.din(w_dff_A_P6cRG2mZ2_0),.clk(gclk));
	jdff dff_A_EMu4TDRX3_0(.dout(w_dff_A_P6cRG2mZ2_0),.din(w_dff_A_EMu4TDRX3_0),.clk(gclk));
	jdff dff_A_AK3xpoD71_0(.dout(w_dff_A_EMu4TDRX3_0),.din(w_dff_A_AK3xpoD71_0),.clk(gclk));
	jdff dff_A_xFjWKTk92_0(.dout(w_dff_A_AK3xpoD71_0),.din(w_dff_A_xFjWKTk92_0),.clk(gclk));
	jdff dff_A_paJVS0G39_0(.dout(w_dff_A_xFjWKTk92_0),.din(w_dff_A_paJVS0G39_0),.clk(gclk));
	jdff dff_A_8VO8diVD1_0(.dout(w_dff_A_paJVS0G39_0),.din(w_dff_A_8VO8diVD1_0),.clk(gclk));
	jdff dff_A_asTtwopN9_0(.dout(w_dff_A_8VO8diVD1_0),.din(w_dff_A_asTtwopN9_0),.clk(gclk));
	jdff dff_B_i2Mv9mSE2_0(.din(n161),.dout(w_dff_B_i2Mv9mSE2_0),.clk(gclk));
	jdff dff_A_7unGc1N81_0(.dout(w_n184_0[0]),.din(w_dff_A_7unGc1N81_0),.clk(gclk));
	jdff dff_A_Ift1tEiP2_0(.dout(w_dff_A_7unGc1N81_0),.din(w_dff_A_Ift1tEiP2_0),.clk(gclk));
	jdff dff_A_WhzBcMHk9_0(.dout(w_dff_A_Ift1tEiP2_0),.din(w_dff_A_WhzBcMHk9_0),.clk(gclk));
	jdff dff_A_QRlEQHcp2_2(.dout(w_n184_0[2]),.din(w_dff_A_QRlEQHcp2_2),.clk(gclk));
	jdff dff_A_fGHsChWy1_2(.dout(w_dff_A_QRlEQHcp2_2),.din(w_dff_A_fGHsChWy1_2),.clk(gclk));
	jdff dff_A_F0a4qMEL1_2(.dout(w_dff_A_fGHsChWy1_2),.din(w_dff_A_F0a4qMEL1_2),.clk(gclk));
	jdff dff_A_USYzVecP0_1(.dout(w_n159_0[1]),.din(w_dff_A_USYzVecP0_1),.clk(gclk));
	jdff dff_A_rIbjrGUp0_0(.dout(w_Gid11_0[0]),.din(w_dff_A_rIbjrGUp0_0),.clk(gclk));
	jdff dff_A_FMIl07QG2_0(.dout(w_dff_A_rIbjrGUp0_0),.din(w_dff_A_FMIl07QG2_0),.clk(gclk));
	jdff dff_A_9OeaZVPh4_0(.dout(w_dff_A_FMIl07QG2_0),.din(w_dff_A_9OeaZVPh4_0),.clk(gclk));
	jdff dff_A_jUt0qhEZ6_0(.dout(w_dff_A_9OeaZVPh4_0),.din(w_dff_A_jUt0qhEZ6_0),.clk(gclk));
	jdff dff_A_HWifq8Fu0_0(.dout(w_dff_A_jUt0qhEZ6_0),.din(w_dff_A_HWifq8Fu0_0),.clk(gclk));
	jdff dff_A_O0Z7EDWG0_0(.dout(w_dff_A_HWifq8Fu0_0),.din(w_dff_A_O0Z7EDWG0_0),.clk(gclk));
	jdff dff_A_9WsiYxJS2_0(.dout(w_dff_A_O0Z7EDWG0_0),.din(w_dff_A_9WsiYxJS2_0),.clk(gclk));
	jdff dff_A_3y2Q2Tqr1_0(.dout(w_dff_A_9WsiYxJS2_0),.din(w_dff_A_3y2Q2Tqr1_0),.clk(gclk));
	jdff dff_A_Lni5NrPW5_0(.dout(w_dff_A_3y2Q2Tqr1_0),.din(w_dff_A_Lni5NrPW5_0),.clk(gclk));
	jdff dff_A_cYKSY5fp6_0(.dout(w_Gid3_0[0]),.din(w_dff_A_cYKSY5fp6_0),.clk(gclk));
	jdff dff_A_ZkJbhuKU3_0(.dout(w_dff_A_cYKSY5fp6_0),.din(w_dff_A_ZkJbhuKU3_0),.clk(gclk));
	jdff dff_A_dRNxF2B02_0(.dout(w_dff_A_ZkJbhuKU3_0),.din(w_dff_A_dRNxF2B02_0),.clk(gclk));
	jdff dff_A_k5Rv8Bkw2_0(.dout(w_dff_A_dRNxF2B02_0),.din(w_dff_A_k5Rv8Bkw2_0),.clk(gclk));
	jdff dff_A_kjRatyLr2_0(.dout(w_dff_A_k5Rv8Bkw2_0),.din(w_dff_A_kjRatyLr2_0),.clk(gclk));
	jdff dff_A_o23deXt75_0(.dout(w_dff_A_kjRatyLr2_0),.din(w_dff_A_o23deXt75_0),.clk(gclk));
	jdff dff_A_L1GO89uh6_0(.dout(w_dff_A_o23deXt75_0),.din(w_dff_A_L1GO89uh6_0),.clk(gclk));
	jdff dff_A_srLF8pSZ3_0(.dout(w_dff_A_L1GO89uh6_0),.din(w_dff_A_srLF8pSZ3_0),.clk(gclk));
	jdff dff_A_jJuM7kdD5_0(.dout(w_dff_A_srLF8pSZ3_0),.din(w_dff_A_jJuM7kdD5_0),.clk(gclk));
	jdff dff_B_nOPe9sMB7_0(.din(n153),.dout(w_dff_B_nOPe9sMB7_0),.clk(gclk));
	jdff dff_B_UC88yyfr6_2(.din(n250),.dout(w_dff_B_UC88yyfr6_2),.clk(gclk));
	jdff dff_A_7GG0Pdeh6_0(.dout(w_n178_0[0]),.din(w_dff_A_7GG0Pdeh6_0),.clk(gclk));
	jdff dff_A_W1UZUwC65_0(.dout(w_dff_A_7GG0Pdeh6_0),.din(w_dff_A_W1UZUwC65_0),.clk(gclk));
	jdff dff_A_d3Pa53nW2_0(.dout(w_dff_A_W1UZUwC65_0),.din(w_dff_A_d3Pa53nW2_0),.clk(gclk));
	jdff dff_A_AaNgmwLP3_2(.dout(w_n178_0[2]),.din(w_dff_A_AaNgmwLP3_2),.clk(gclk));
	jdff dff_A_8iiCmORe1_2(.dout(w_dff_A_AaNgmwLP3_2),.din(w_dff_A_8iiCmORe1_2),.clk(gclk));
	jdff dff_A_vdMCMSdo5_2(.dout(w_dff_A_8iiCmORe1_2),.din(w_dff_A_vdMCMSdo5_2),.clk(gclk));
	jdff dff_A_7VTeUlZZ6_1(.dout(w_n150_0[1]),.din(w_dff_A_7VTeUlZZ6_1),.clk(gclk));
	jdff dff_A_eIv5XzI46_0(.dout(w_Gid9_0[0]),.din(w_dff_A_eIv5XzI46_0),.clk(gclk));
	jdff dff_A_O76DOFuz5_0(.dout(w_dff_A_eIv5XzI46_0),.din(w_dff_A_O76DOFuz5_0),.clk(gclk));
	jdff dff_A_A4go7Xc77_0(.dout(w_dff_A_O76DOFuz5_0),.din(w_dff_A_A4go7Xc77_0),.clk(gclk));
	jdff dff_A_6NZCI8ZK6_0(.dout(w_dff_A_A4go7Xc77_0),.din(w_dff_A_6NZCI8ZK6_0),.clk(gclk));
	jdff dff_A_j2adSQB68_0(.dout(w_dff_A_6NZCI8ZK6_0),.din(w_dff_A_j2adSQB68_0),.clk(gclk));
	jdff dff_A_djVnZcu11_0(.dout(w_dff_A_j2adSQB68_0),.din(w_dff_A_djVnZcu11_0),.clk(gclk));
	jdff dff_A_Ug0wiIoZ7_0(.dout(w_dff_A_djVnZcu11_0),.din(w_dff_A_Ug0wiIoZ7_0),.clk(gclk));
	jdff dff_A_3lXIVw5j2_0(.dout(w_dff_A_Ug0wiIoZ7_0),.din(w_dff_A_3lXIVw5j2_0),.clk(gclk));
	jdff dff_A_KnxHH5LI4_0(.dout(w_dff_A_3lXIVw5j2_0),.din(w_dff_A_KnxHH5LI4_0),.clk(gclk));
	jdff dff_A_1dR3VcGE8_0(.dout(w_Gid1_0[0]),.din(w_dff_A_1dR3VcGE8_0),.clk(gclk));
	jdff dff_A_PLZhoxte0_0(.dout(w_dff_A_1dR3VcGE8_0),.din(w_dff_A_PLZhoxte0_0),.clk(gclk));
	jdff dff_A_tlO5yp5z1_0(.dout(w_dff_A_PLZhoxte0_0),.din(w_dff_A_tlO5yp5z1_0),.clk(gclk));
	jdff dff_A_gSm9D3Ag9_0(.dout(w_dff_A_tlO5yp5z1_0),.din(w_dff_A_gSm9D3Ag9_0),.clk(gclk));
	jdff dff_A_Sq4JzbZU8_0(.dout(w_dff_A_gSm9D3Ag9_0),.din(w_dff_A_Sq4JzbZU8_0),.clk(gclk));
	jdff dff_A_V7qKu6Bj9_0(.dout(w_dff_A_Sq4JzbZU8_0),.din(w_dff_A_V7qKu6Bj9_0),.clk(gclk));
	jdff dff_A_PyxwTlgq3_0(.dout(w_dff_A_V7qKu6Bj9_0),.din(w_dff_A_PyxwTlgq3_0),.clk(gclk));
	jdff dff_A_eZFHzSBZ1_0(.dout(w_dff_A_PyxwTlgq3_0),.din(w_dff_A_eZFHzSBZ1_0),.clk(gclk));
	jdff dff_A_ibDwxNCx3_0(.dout(w_dff_A_eZFHzSBZ1_0),.din(w_dff_A_ibDwxNCx3_0),.clk(gclk));
	jdff dff_A_lxrLuyYV2_0(.dout(w_Gid26_0[0]),.din(w_dff_A_lxrLuyYV2_0),.clk(gclk));
	jdff dff_A_HaVaPBOT7_0(.dout(w_dff_A_lxrLuyYV2_0),.din(w_dff_A_HaVaPBOT7_0),.clk(gclk));
	jdff dff_A_MbULmuV91_0(.dout(w_dff_A_HaVaPBOT7_0),.din(w_dff_A_MbULmuV91_0),.clk(gclk));
	jdff dff_A_FCbjU2kj8_0(.dout(w_dff_A_MbULmuV91_0),.din(w_dff_A_FCbjU2kj8_0),.clk(gclk));
	jdff dff_A_y728LCBF3_0(.dout(w_dff_A_FCbjU2kj8_0),.din(w_dff_A_y728LCBF3_0),.clk(gclk));
	jdff dff_A_wRXh8FI02_0(.dout(w_dff_A_y728LCBF3_0),.din(w_dff_A_wRXh8FI02_0),.clk(gclk));
	jdff dff_A_4tyfHfTH3_0(.dout(w_dff_A_wRXh8FI02_0),.din(w_dff_A_4tyfHfTH3_0),.clk(gclk));
	jdff dff_A_RflG3I773_0(.dout(w_dff_A_4tyfHfTH3_0),.din(w_dff_A_RflG3I773_0),.clk(gclk));
	jdff dff_A_mLEMYJRM9_0(.dout(w_dff_A_RflG3I773_0),.din(w_dff_A_mLEMYJRM9_0),.clk(gclk));
	jdff dff_A_MRxFezn76_0(.dout(w_Gid25_0[0]),.din(w_dff_A_MRxFezn76_0),.clk(gclk));
	jdff dff_A_AnF5QnyT9_0(.dout(w_dff_A_MRxFezn76_0),.din(w_dff_A_AnF5QnyT9_0),.clk(gclk));
	jdff dff_A_pxK0fo0l9_0(.dout(w_dff_A_AnF5QnyT9_0),.din(w_dff_A_pxK0fo0l9_0),.clk(gclk));
	jdff dff_A_slVlHIJ22_0(.dout(w_dff_A_pxK0fo0l9_0),.din(w_dff_A_slVlHIJ22_0),.clk(gclk));
	jdff dff_A_UhdG2aDJ3_0(.dout(w_dff_A_slVlHIJ22_0),.din(w_dff_A_UhdG2aDJ3_0),.clk(gclk));
	jdff dff_A_qf8HLpB87_0(.dout(w_dff_A_UhdG2aDJ3_0),.din(w_dff_A_qf8HLpB87_0),.clk(gclk));
	jdff dff_A_hk1hBb262_0(.dout(w_dff_A_qf8HLpB87_0),.din(w_dff_A_hk1hBb262_0),.clk(gclk));
	jdff dff_A_s3aYkSp83_0(.dout(w_dff_A_hk1hBb262_0),.din(w_dff_A_s3aYkSp83_0),.clk(gclk));
	jdff dff_A_p0JsYRz87_0(.dout(w_dff_A_s3aYkSp83_0),.din(w_dff_A_p0JsYRz87_0),.clk(gclk));
	jdff dff_A_lD0vxeIb6_0(.dout(w_Gid24_0[0]),.din(w_dff_A_lD0vxeIb6_0),.clk(gclk));
	jdff dff_A_zVPlDPcz1_0(.dout(w_dff_A_lD0vxeIb6_0),.din(w_dff_A_zVPlDPcz1_0),.clk(gclk));
	jdff dff_A_Szl2p8Dp3_0(.dout(w_dff_A_zVPlDPcz1_0),.din(w_dff_A_Szl2p8Dp3_0),.clk(gclk));
	jdff dff_A_y2fbIcPa9_0(.dout(w_dff_A_Szl2p8Dp3_0),.din(w_dff_A_y2fbIcPa9_0),.clk(gclk));
	jdff dff_A_ZIWQSUWm1_0(.dout(w_dff_A_y2fbIcPa9_0),.din(w_dff_A_ZIWQSUWm1_0),.clk(gclk));
	jdff dff_A_0mxIEL0Z9_0(.dout(w_dff_A_ZIWQSUWm1_0),.din(w_dff_A_0mxIEL0Z9_0),.clk(gclk));
	jdff dff_A_ZeTrkn1Q2_0(.dout(w_dff_A_0mxIEL0Z9_0),.din(w_dff_A_ZeTrkn1Q2_0),.clk(gclk));
	jdff dff_A_kdFYze5e1_0(.dout(w_dff_A_ZeTrkn1Q2_0),.din(w_dff_A_kdFYze5e1_0),.clk(gclk));
	jdff dff_A_2bZYM1jj9_0(.dout(w_dff_A_kdFYze5e1_0),.din(w_dff_A_2bZYM1jj9_0),.clk(gclk));
	jdff dff_B_fq2pqfIy1_1(.din(n138),.dout(w_dff_B_fq2pqfIy1_1),.clk(gclk));
	jdff dff_A_PrT5yRJK7_0(.dout(w_Gid30_0[0]),.din(w_dff_A_PrT5yRJK7_0),.clk(gclk));
	jdff dff_A_K4S6b3Qc3_0(.dout(w_dff_A_PrT5yRJK7_0),.din(w_dff_A_K4S6b3Qc3_0),.clk(gclk));
	jdff dff_A_oPbRgCbe7_0(.dout(w_dff_A_K4S6b3Qc3_0),.din(w_dff_A_oPbRgCbe7_0),.clk(gclk));
	jdff dff_A_6k88Ow9F8_0(.dout(w_dff_A_oPbRgCbe7_0),.din(w_dff_A_6k88Ow9F8_0),.clk(gclk));
	jdff dff_A_JJJrjD4X6_0(.dout(w_dff_A_6k88Ow9F8_0),.din(w_dff_A_JJJrjD4X6_0),.clk(gclk));
	jdff dff_A_4iWHi9c62_0(.dout(w_dff_A_JJJrjD4X6_0),.din(w_dff_A_4iWHi9c62_0),.clk(gclk));
	jdff dff_A_JmYSlVj16_0(.dout(w_dff_A_4iWHi9c62_0),.din(w_dff_A_JmYSlVj16_0),.clk(gclk));
	jdff dff_A_9f7E5E7Q2_0(.dout(w_dff_A_JmYSlVj16_0),.din(w_dff_A_9f7E5E7Q2_0),.clk(gclk));
	jdff dff_A_PGuNR5kM5_0(.dout(w_dff_A_9f7E5E7Q2_0),.din(w_dff_A_PGuNR5kM5_0),.clk(gclk));
	jdff dff_A_Ks24DUMm1_0(.dout(w_Gid29_0[0]),.din(w_dff_A_Ks24DUMm1_0),.clk(gclk));
	jdff dff_A_2b1dVPwE6_0(.dout(w_dff_A_Ks24DUMm1_0),.din(w_dff_A_2b1dVPwE6_0),.clk(gclk));
	jdff dff_A_OR7hYgjl6_0(.dout(w_dff_A_2b1dVPwE6_0),.din(w_dff_A_OR7hYgjl6_0),.clk(gclk));
	jdff dff_A_dn89tSFB9_0(.dout(w_dff_A_OR7hYgjl6_0),.din(w_dff_A_dn89tSFB9_0),.clk(gclk));
	jdff dff_A_A0n2jZf65_0(.dout(w_dff_A_dn89tSFB9_0),.din(w_dff_A_A0n2jZf65_0),.clk(gclk));
	jdff dff_A_EqzUeRIk8_0(.dout(w_dff_A_A0n2jZf65_0),.din(w_dff_A_EqzUeRIk8_0),.clk(gclk));
	jdff dff_A_Uj4GsI588_0(.dout(w_dff_A_EqzUeRIk8_0),.din(w_dff_A_Uj4GsI588_0),.clk(gclk));
	jdff dff_A_LWVePi6g3_0(.dout(w_dff_A_Uj4GsI588_0),.din(w_dff_A_LWVePi6g3_0),.clk(gclk));
	jdff dff_A_lpdSTX472_0(.dout(w_dff_A_LWVePi6g3_0),.din(w_dff_A_lpdSTX472_0),.clk(gclk));
	jdff dff_A_x2JCpfEA2_0(.dout(w_Gid28_0[0]),.din(w_dff_A_x2JCpfEA2_0),.clk(gclk));
	jdff dff_A_CRzMu6Ej3_0(.dout(w_dff_A_x2JCpfEA2_0),.din(w_dff_A_CRzMu6Ej3_0),.clk(gclk));
	jdff dff_A_t0ciBwgo1_0(.dout(w_dff_A_CRzMu6Ej3_0),.din(w_dff_A_t0ciBwgo1_0),.clk(gclk));
	jdff dff_A_HgWc9BkZ2_0(.dout(w_dff_A_t0ciBwgo1_0),.din(w_dff_A_HgWc9BkZ2_0),.clk(gclk));
	jdff dff_A_KIJqRfKM4_0(.dout(w_dff_A_HgWc9BkZ2_0),.din(w_dff_A_KIJqRfKM4_0),.clk(gclk));
	jdff dff_A_2vN6qVH66_0(.dout(w_dff_A_KIJqRfKM4_0),.din(w_dff_A_2vN6qVH66_0),.clk(gclk));
	jdff dff_A_tavcwFC29_0(.dout(w_dff_A_2vN6qVH66_0),.din(w_dff_A_tavcwFC29_0),.clk(gclk));
	jdff dff_A_ALXC0HG02_0(.dout(w_dff_A_tavcwFC29_0),.din(w_dff_A_ALXC0HG02_0),.clk(gclk));
	jdff dff_A_KqvraJus8_0(.dout(w_dff_A_ALXC0HG02_0),.din(w_dff_A_KqvraJus8_0),.clk(gclk));
	jdff dff_A_PXTVRGeM9_1(.dout(w_n87_0[1]),.din(w_dff_A_PXTVRGeM9_1),.clk(gclk));
	jdff dff_A_1FxENjWr2_0(.dout(w_Gid22_0[0]),.din(w_dff_A_1FxENjWr2_0),.clk(gclk));
	jdff dff_A_ogf2vX5S4_0(.dout(w_dff_A_1FxENjWr2_0),.din(w_dff_A_ogf2vX5S4_0),.clk(gclk));
	jdff dff_A_jqihCHYU0_0(.dout(w_dff_A_ogf2vX5S4_0),.din(w_dff_A_jqihCHYU0_0),.clk(gclk));
	jdff dff_A_T0SHlAxV4_0(.dout(w_dff_A_jqihCHYU0_0),.din(w_dff_A_T0SHlAxV4_0),.clk(gclk));
	jdff dff_A_WFMAe56z7_0(.dout(w_dff_A_T0SHlAxV4_0),.din(w_dff_A_WFMAe56z7_0),.clk(gclk));
	jdff dff_A_kTa85LaC5_0(.dout(w_dff_A_WFMAe56z7_0),.din(w_dff_A_kTa85LaC5_0),.clk(gclk));
	jdff dff_A_uvTLUANg3_0(.dout(w_dff_A_kTa85LaC5_0),.din(w_dff_A_uvTLUANg3_0),.clk(gclk));
	jdff dff_A_gZbEjkNZ1_0(.dout(w_dff_A_uvTLUANg3_0),.din(w_dff_A_gZbEjkNZ1_0),.clk(gclk));
	jdff dff_A_ZlF6DRNS8_0(.dout(w_dff_A_gZbEjkNZ1_0),.din(w_dff_A_ZlF6DRNS8_0),.clk(gclk));
	jdff dff_A_tiBLV1YL1_0(.dout(w_Gid21_0[0]),.din(w_dff_A_tiBLV1YL1_0),.clk(gclk));
	jdff dff_A_1rqcKS623_0(.dout(w_dff_A_tiBLV1YL1_0),.din(w_dff_A_1rqcKS623_0),.clk(gclk));
	jdff dff_A_FovqzTDo5_0(.dout(w_dff_A_1rqcKS623_0),.din(w_dff_A_FovqzTDo5_0),.clk(gclk));
	jdff dff_A_ObNp9zp69_0(.dout(w_dff_A_FovqzTDo5_0),.din(w_dff_A_ObNp9zp69_0),.clk(gclk));
	jdff dff_A_YJG9NDrE3_0(.dout(w_dff_A_ObNp9zp69_0),.din(w_dff_A_YJG9NDrE3_0),.clk(gclk));
	jdff dff_A_Zwo4CKf33_0(.dout(w_dff_A_YJG9NDrE3_0),.din(w_dff_A_Zwo4CKf33_0),.clk(gclk));
	jdff dff_A_rx7JAJlH8_0(.dout(w_dff_A_Zwo4CKf33_0),.din(w_dff_A_rx7JAJlH8_0),.clk(gclk));
	jdff dff_A_nhJEgkeJ4_0(.dout(w_dff_A_rx7JAJlH8_0),.din(w_dff_A_nhJEgkeJ4_0),.clk(gclk));
	jdff dff_A_SBxBORC27_0(.dout(w_dff_A_nhJEgkeJ4_0),.din(w_dff_A_SBxBORC27_0),.clk(gclk));
	jdff dff_A_tV8yo2h87_0(.dout(w_Gid20_0[0]),.din(w_dff_A_tV8yo2h87_0),.clk(gclk));
	jdff dff_A_buwdRfLs2_0(.dout(w_dff_A_tV8yo2h87_0),.din(w_dff_A_buwdRfLs2_0),.clk(gclk));
	jdff dff_A_B0zqrSuL5_0(.dout(w_dff_A_buwdRfLs2_0),.din(w_dff_A_B0zqrSuL5_0),.clk(gclk));
	jdff dff_A_eiyFXXyB3_0(.dout(w_dff_A_B0zqrSuL5_0),.din(w_dff_A_eiyFXXyB3_0),.clk(gclk));
	jdff dff_A_AggnXpA57_0(.dout(w_dff_A_eiyFXXyB3_0),.din(w_dff_A_AggnXpA57_0),.clk(gclk));
	jdff dff_A_t9LVRxAo2_0(.dout(w_dff_A_AggnXpA57_0),.din(w_dff_A_t9LVRxAo2_0),.clk(gclk));
	jdff dff_A_EhC0h2vs5_0(.dout(w_dff_A_t9LVRxAo2_0),.din(w_dff_A_EhC0h2vs5_0),.clk(gclk));
	jdff dff_A_j0D5SOUx4_0(.dout(w_dff_A_EhC0h2vs5_0),.din(w_dff_A_j0D5SOUx4_0),.clk(gclk));
	jdff dff_A_8AF4rwWG4_0(.dout(w_dff_A_j0D5SOUx4_0),.din(w_dff_A_8AF4rwWG4_0),.clk(gclk));
	jdff dff_A_0IZLWlvP1_0(.dout(w_Gid8_0[0]),.din(w_dff_A_0IZLWlvP1_0),.clk(gclk));
	jdff dff_A_B860Ugzw7_0(.dout(w_dff_A_0IZLWlvP1_0),.din(w_dff_A_B860Ugzw7_0),.clk(gclk));
	jdff dff_A_zgh7f9YY9_0(.dout(w_dff_A_B860Ugzw7_0),.din(w_dff_A_zgh7f9YY9_0),.clk(gclk));
	jdff dff_A_GoHujcHd9_0(.dout(w_dff_A_zgh7f9YY9_0),.din(w_dff_A_GoHujcHd9_0),.clk(gclk));
	jdff dff_A_GoZClivP6_0(.dout(w_dff_A_GoHujcHd9_0),.din(w_dff_A_GoZClivP6_0),.clk(gclk));
	jdff dff_A_S8VSJANp4_0(.dout(w_dff_A_GoZClivP6_0),.din(w_dff_A_S8VSJANp4_0),.clk(gclk));
	jdff dff_A_6YWNRBmi0_0(.dout(w_dff_A_S8VSJANp4_0),.din(w_dff_A_6YWNRBmi0_0),.clk(gclk));
	jdff dff_A_Mo7Czp4I5_0(.dout(w_dff_A_6YWNRBmi0_0),.din(w_dff_A_Mo7Czp4I5_0),.clk(gclk));
	jdff dff_A_Fm81bVXb4_0(.dout(w_dff_A_Mo7Czp4I5_0),.din(w_dff_A_Fm81bVXb4_0),.clk(gclk));
	jdff dff_A_rTsSmuLl0_0(.dout(w_Gid0_0[0]),.din(w_dff_A_rTsSmuLl0_0),.clk(gclk));
	jdff dff_A_5BQ3PXpO5_0(.dout(w_dff_A_rTsSmuLl0_0),.din(w_dff_A_5BQ3PXpO5_0),.clk(gclk));
	jdff dff_A_WTIBzFbc1_0(.dout(w_dff_A_5BQ3PXpO5_0),.din(w_dff_A_WTIBzFbc1_0),.clk(gclk));
	jdff dff_A_0JzMntPC8_0(.dout(w_dff_A_WTIBzFbc1_0),.din(w_dff_A_0JzMntPC8_0),.clk(gclk));
	jdff dff_A_NogwJga58_0(.dout(w_dff_A_0JzMntPC8_0),.din(w_dff_A_NogwJga58_0),.clk(gclk));
	jdff dff_A_6pFiOnxD8_0(.dout(w_dff_A_NogwJga58_0),.din(w_dff_A_6pFiOnxD8_0),.clk(gclk));
	jdff dff_A_eMP34gdl6_0(.dout(w_dff_A_6pFiOnxD8_0),.din(w_dff_A_eMP34gdl6_0),.clk(gclk));
	jdff dff_A_vFmJqvz96_0(.dout(w_dff_A_eMP34gdl6_0),.din(w_dff_A_vFmJqvz96_0),.clk(gclk));
	jdff dff_A_jeIqdny36_0(.dout(w_dff_A_vFmJqvz96_0),.din(w_dff_A_jeIqdny36_0),.clk(gclk));
	jdff dff_B_cIPsQN239_1(.din(n75),.dout(w_dff_B_cIPsQN239_1),.clk(gclk));
	jdff dff_A_LWCSZxky9_0(.dout(w_Gid18_0[0]),.din(w_dff_A_LWCSZxky9_0),.clk(gclk));
	jdff dff_A_CtBCDOTn2_0(.dout(w_dff_A_LWCSZxky9_0),.din(w_dff_A_CtBCDOTn2_0),.clk(gclk));
	jdff dff_A_0AKNiRU74_0(.dout(w_dff_A_CtBCDOTn2_0),.din(w_dff_A_0AKNiRU74_0),.clk(gclk));
	jdff dff_A_r4oiOSDq0_0(.dout(w_dff_A_0AKNiRU74_0),.din(w_dff_A_r4oiOSDq0_0),.clk(gclk));
	jdff dff_A_YDvw6Okc5_0(.dout(w_dff_A_r4oiOSDq0_0),.din(w_dff_A_YDvw6Okc5_0),.clk(gclk));
	jdff dff_A_yjVHrI783_0(.dout(w_dff_A_YDvw6Okc5_0),.din(w_dff_A_yjVHrI783_0),.clk(gclk));
	jdff dff_A_8aYyWgMp2_0(.dout(w_dff_A_yjVHrI783_0),.din(w_dff_A_8aYyWgMp2_0),.clk(gclk));
	jdff dff_A_hyVhuwv11_0(.dout(w_dff_A_8aYyWgMp2_0),.din(w_dff_A_hyVhuwv11_0),.clk(gclk));
	jdff dff_A_pEGxduJo7_0(.dout(w_dff_A_hyVhuwv11_0),.din(w_dff_A_pEGxduJo7_0),.clk(gclk));
	jdff dff_A_YtPkck9X0_0(.dout(w_Gid17_0[0]),.din(w_dff_A_YtPkck9X0_0),.clk(gclk));
	jdff dff_A_3GW6Q84W5_0(.dout(w_dff_A_YtPkck9X0_0),.din(w_dff_A_3GW6Q84W5_0),.clk(gclk));
	jdff dff_A_xlCckJXS9_0(.dout(w_dff_A_3GW6Q84W5_0),.din(w_dff_A_xlCckJXS9_0),.clk(gclk));
	jdff dff_A_Eqxn9ihg9_0(.dout(w_dff_A_xlCckJXS9_0),.din(w_dff_A_Eqxn9ihg9_0),.clk(gclk));
	jdff dff_A_09sQ4T991_0(.dout(w_dff_A_Eqxn9ihg9_0),.din(w_dff_A_09sQ4T991_0),.clk(gclk));
	jdff dff_A_jinmfTAn7_0(.dout(w_dff_A_09sQ4T991_0),.din(w_dff_A_jinmfTAn7_0),.clk(gclk));
	jdff dff_A_tIx9bA3Q0_0(.dout(w_dff_A_jinmfTAn7_0),.din(w_dff_A_tIx9bA3Q0_0),.clk(gclk));
	jdff dff_A_w8A5x5PP4_0(.dout(w_dff_A_tIx9bA3Q0_0),.din(w_dff_A_w8A5x5PP4_0),.clk(gclk));
	jdff dff_A_TLDVzjjS5_0(.dout(w_dff_A_w8A5x5PP4_0),.din(w_dff_A_TLDVzjjS5_0),.clk(gclk));
	jdff dff_A_Pm24qRSh2_0(.dout(w_Gid16_0[0]),.din(w_dff_A_Pm24qRSh2_0),.clk(gclk));
	jdff dff_A_UQ6moDOL1_0(.dout(w_dff_A_Pm24qRSh2_0),.din(w_dff_A_UQ6moDOL1_0),.clk(gclk));
	jdff dff_A_DunxYemY2_0(.dout(w_dff_A_UQ6moDOL1_0),.din(w_dff_A_DunxYemY2_0),.clk(gclk));
	jdff dff_A_2aI3FGae6_0(.dout(w_dff_A_DunxYemY2_0),.din(w_dff_A_2aI3FGae6_0),.clk(gclk));
	jdff dff_A_IsXqFmFF4_0(.dout(w_dff_A_2aI3FGae6_0),.din(w_dff_A_IsXqFmFF4_0),.clk(gclk));
	jdff dff_A_561XGa8Q4_0(.dout(w_dff_A_IsXqFmFF4_0),.din(w_dff_A_561XGa8Q4_0),.clk(gclk));
	jdff dff_A_XfgkVAcc8_0(.dout(w_dff_A_561XGa8Q4_0),.din(w_dff_A_XfgkVAcc8_0),.clk(gclk));
	jdff dff_A_c6GpQIdt8_0(.dout(w_dff_A_XfgkVAcc8_0),.din(w_dff_A_c6GpQIdt8_0),.clk(gclk));
	jdff dff_A_7a90pXgD9_0(.dout(w_dff_A_c6GpQIdt8_0),.din(w_dff_A_7a90pXgD9_0),.clk(gclk));
	jdff dff_A_k0bCiLaS2_1(.dout(w_n187_0[1]),.din(w_dff_A_k0bCiLaS2_1),.clk(gclk));
	jdff dff_A_f2s8mWow7_1(.dout(w_dff_A_k0bCiLaS2_1),.din(w_dff_A_f2s8mWow7_1),.clk(gclk));
	jdff dff_A_5g65sS2q0_1(.dout(w_dff_A_f2s8mWow7_1),.din(w_dff_A_5g65sS2q0_1),.clk(gclk));
	jdff dff_A_kCJ787kt9_2(.dout(w_n187_0[2]),.din(w_dff_A_kCJ787kt9_2),.clk(gclk));
	jdff dff_A_8aSTICIo0_2(.dout(w_dff_A_kCJ787kt9_2),.din(w_dff_A_8aSTICIo0_2),.clk(gclk));
	jdff dff_A_SI7LRVvI5_2(.dout(w_dff_A_8aSTICIo0_2),.din(w_dff_A_SI7LRVvI5_2),.clk(gclk));
	jdff dff_A_onFBGz5h5_1(.dout(w_n102_1[1]),.din(w_dff_A_onFBGz5h5_1),.clk(gclk));
	jdff dff_A_ahfjs8qw3_0(.dout(w_Gid31_0[0]),.din(w_dff_A_ahfjs8qw3_0),.clk(gclk));
	jdff dff_A_4CBE20Fx6_0(.dout(w_dff_A_ahfjs8qw3_0),.din(w_dff_A_4CBE20Fx6_0),.clk(gclk));
	jdff dff_A_CmfBq9W25_0(.dout(w_dff_A_4CBE20Fx6_0),.din(w_dff_A_CmfBq9W25_0),.clk(gclk));
	jdff dff_A_VkDfYNUq3_0(.dout(w_dff_A_CmfBq9W25_0),.din(w_dff_A_VkDfYNUq3_0),.clk(gclk));
	jdff dff_A_986HQcMu7_0(.dout(w_dff_A_VkDfYNUq3_0),.din(w_dff_A_986HQcMu7_0),.clk(gclk));
	jdff dff_A_7atJrpkP6_0(.dout(w_dff_A_986HQcMu7_0),.din(w_dff_A_7atJrpkP6_0),.clk(gclk));
	jdff dff_A_wIzZywLv4_0(.dout(w_dff_A_7atJrpkP6_0),.din(w_dff_A_wIzZywLv4_0),.clk(gclk));
	jdff dff_A_2n5YP8lt9_0(.dout(w_dff_A_wIzZywLv4_0),.din(w_dff_A_2n5YP8lt9_0),.clk(gclk));
	jdff dff_A_Mk7fOtus9_0(.dout(w_dff_A_2n5YP8lt9_0),.din(w_dff_A_Mk7fOtus9_0),.clk(gclk));
	jdff dff_A_Iobxln0X2_0(.dout(w_Gid27_0[0]),.din(w_dff_A_Iobxln0X2_0),.clk(gclk));
	jdff dff_A_y74magwy5_0(.dout(w_dff_A_Iobxln0X2_0),.din(w_dff_A_y74magwy5_0),.clk(gclk));
	jdff dff_A_EBxyZdkC6_0(.dout(w_dff_A_y74magwy5_0),.din(w_dff_A_EBxyZdkC6_0),.clk(gclk));
	jdff dff_A_4WUkd2ps2_0(.dout(w_dff_A_EBxyZdkC6_0),.din(w_dff_A_4WUkd2ps2_0),.clk(gclk));
	jdff dff_A_glBX3B5F6_0(.dout(w_dff_A_4WUkd2ps2_0),.din(w_dff_A_glBX3B5F6_0),.clk(gclk));
	jdff dff_A_aYEnnFAd7_0(.dout(w_dff_A_glBX3B5F6_0),.din(w_dff_A_aYEnnFAd7_0),.clk(gclk));
	jdff dff_A_k6sA7Hxe1_0(.dout(w_dff_A_aYEnnFAd7_0),.din(w_dff_A_k6sA7Hxe1_0),.clk(gclk));
	jdff dff_A_yhkskwpx8_0(.dout(w_dff_A_k6sA7Hxe1_0),.din(w_dff_A_yhkskwpx8_0),.clk(gclk));
	jdff dff_A_atPkpVhr5_0(.dout(w_dff_A_yhkskwpx8_0),.din(w_dff_A_atPkpVhr5_0),.clk(gclk));
	jdff dff_A_xQ0AQxpe6_0(.dout(w_Gid23_0[0]),.din(w_dff_A_xQ0AQxpe6_0),.clk(gclk));
	jdff dff_A_9X4gwM5a4_0(.dout(w_dff_A_xQ0AQxpe6_0),.din(w_dff_A_9X4gwM5a4_0),.clk(gclk));
	jdff dff_A_lo9aW5vm6_0(.dout(w_dff_A_9X4gwM5a4_0),.din(w_dff_A_lo9aW5vm6_0),.clk(gclk));
	jdff dff_A_IVsM3AX00_0(.dout(w_dff_A_lo9aW5vm6_0),.din(w_dff_A_IVsM3AX00_0),.clk(gclk));
	jdff dff_A_7WgGb0fo2_0(.dout(w_dff_A_IVsM3AX00_0),.din(w_dff_A_7WgGb0fo2_0),.clk(gclk));
	jdff dff_A_v6WQ1kX65_0(.dout(w_dff_A_7WgGb0fo2_0),.din(w_dff_A_v6WQ1kX65_0),.clk(gclk));
	jdff dff_A_NDLb4voV1_0(.dout(w_dff_A_v6WQ1kX65_0),.din(w_dff_A_NDLb4voV1_0),.clk(gclk));
	jdff dff_A_pXkblSMP7_0(.dout(w_dff_A_NDLb4voV1_0),.din(w_dff_A_pXkblSMP7_0),.clk(gclk));
	jdff dff_A_PiQJmDTh0_0(.dout(w_dff_A_pXkblSMP7_0),.din(w_dff_A_PiQJmDTh0_0),.clk(gclk));
	jdff dff_A_Q4CMYELA8_0(.dout(w_Gid19_0[0]),.din(w_dff_A_Q4CMYELA8_0),.clk(gclk));
	jdff dff_A_3YawHl5y3_0(.dout(w_dff_A_Q4CMYELA8_0),.din(w_dff_A_3YawHl5y3_0),.clk(gclk));
	jdff dff_A_OKVBf5Ep3_0(.dout(w_dff_A_3YawHl5y3_0),.din(w_dff_A_OKVBf5Ep3_0),.clk(gclk));
	jdff dff_A_vqbeihJG0_0(.dout(w_dff_A_OKVBf5Ep3_0),.din(w_dff_A_vqbeihJG0_0),.clk(gclk));
	jdff dff_A_7rrmaD3S8_0(.dout(w_dff_A_vqbeihJG0_0),.din(w_dff_A_7rrmaD3S8_0),.clk(gclk));
	jdff dff_A_aSyoe34x4_0(.dout(w_dff_A_7rrmaD3S8_0),.din(w_dff_A_aSyoe34x4_0),.clk(gclk));
	jdff dff_A_ooiB0p4j7_0(.dout(w_dff_A_aSyoe34x4_0),.din(w_dff_A_ooiB0p4j7_0),.clk(gclk));
	jdff dff_A_z4c8E6dp7_0(.dout(w_dff_A_ooiB0p4j7_0),.din(w_dff_A_z4c8E6dp7_0),.clk(gclk));
	jdff dff_A_nCnJAGQY6_0(.dout(w_dff_A_z4c8E6dp7_0),.din(w_dff_A_nCnJAGQY6_0),.clk(gclk));
	jdff dff_A_XpIpBYFo4_0(.dout(w_Gid15_0[0]),.din(w_dff_A_XpIpBYFo4_0),.clk(gclk));
	jdff dff_A_SjxrMhjv6_0(.dout(w_dff_A_XpIpBYFo4_0),.din(w_dff_A_SjxrMhjv6_0),.clk(gclk));
	jdff dff_A_diQhLNkK8_0(.dout(w_dff_A_SjxrMhjv6_0),.din(w_dff_A_diQhLNkK8_0),.clk(gclk));
	jdff dff_A_vLDnubxj3_0(.dout(w_dff_A_diQhLNkK8_0),.din(w_dff_A_vLDnubxj3_0),.clk(gclk));
	jdff dff_A_DNmO7cE60_0(.dout(w_dff_A_vLDnubxj3_0),.din(w_dff_A_DNmO7cE60_0),.clk(gclk));
	jdff dff_A_lXkyjtLR9_0(.dout(w_dff_A_DNmO7cE60_0),.din(w_dff_A_lXkyjtLR9_0),.clk(gclk));
	jdff dff_A_dOzgrWnE1_0(.dout(w_dff_A_lXkyjtLR9_0),.din(w_dff_A_dOzgrWnE1_0),.clk(gclk));
	jdff dff_A_0eJjrkoH9_0(.dout(w_dff_A_dOzgrWnE1_0),.din(w_dff_A_0eJjrkoH9_0),.clk(gclk));
	jdff dff_A_4KrvNnKl3_0(.dout(w_dff_A_0eJjrkoH9_0),.din(w_dff_A_4KrvNnKl3_0),.clk(gclk));
	jdff dff_A_6wLaNSOi9_0(.dout(w_Gid14_0[0]),.din(w_dff_A_6wLaNSOi9_0),.clk(gclk));
	jdff dff_A_2kyX6NGj2_0(.dout(w_dff_A_6wLaNSOi9_0),.din(w_dff_A_2kyX6NGj2_0),.clk(gclk));
	jdff dff_A_tGScyidT4_0(.dout(w_dff_A_2kyX6NGj2_0),.din(w_dff_A_tGScyidT4_0),.clk(gclk));
	jdff dff_A_fSged4Wv5_0(.dout(w_dff_A_tGScyidT4_0),.din(w_dff_A_fSged4Wv5_0),.clk(gclk));
	jdff dff_A_Zi3qTDkl0_0(.dout(w_dff_A_fSged4Wv5_0),.din(w_dff_A_Zi3qTDkl0_0),.clk(gclk));
	jdff dff_A_QurSle926_0(.dout(w_dff_A_Zi3qTDkl0_0),.din(w_dff_A_QurSle926_0),.clk(gclk));
	jdff dff_A_3LAcBKPj4_0(.dout(w_dff_A_QurSle926_0),.din(w_dff_A_3LAcBKPj4_0),.clk(gclk));
	jdff dff_A_4GZxTSrF7_0(.dout(w_dff_A_3LAcBKPj4_0),.din(w_dff_A_4GZxTSrF7_0),.clk(gclk));
	jdff dff_A_QIjOxqaN9_0(.dout(w_dff_A_4GZxTSrF7_0),.din(w_dff_A_QIjOxqaN9_0),.clk(gclk));
	jdff dff_A_vh1jU26g1_0(.dout(w_Gid13_0[0]),.din(w_dff_A_vh1jU26g1_0),.clk(gclk));
	jdff dff_A_q1lzO1Xl8_0(.dout(w_dff_A_vh1jU26g1_0),.din(w_dff_A_q1lzO1Xl8_0),.clk(gclk));
	jdff dff_A_MEyKYcYZ2_0(.dout(w_dff_A_q1lzO1Xl8_0),.din(w_dff_A_MEyKYcYZ2_0),.clk(gclk));
	jdff dff_A_GSX6na7u8_0(.dout(w_dff_A_MEyKYcYZ2_0),.din(w_dff_A_GSX6na7u8_0),.clk(gclk));
	jdff dff_A_2o412wT18_0(.dout(w_dff_A_GSX6na7u8_0),.din(w_dff_A_2o412wT18_0),.clk(gclk));
	jdff dff_A_C9yWhCjS6_0(.dout(w_dff_A_2o412wT18_0),.din(w_dff_A_C9yWhCjS6_0),.clk(gclk));
	jdff dff_A_BeOAonQr0_0(.dout(w_dff_A_C9yWhCjS6_0),.din(w_dff_A_BeOAonQr0_0),.clk(gclk));
	jdff dff_A_Vhb6DImv1_0(.dout(w_dff_A_BeOAonQr0_0),.din(w_dff_A_Vhb6DImv1_0),.clk(gclk));
	jdff dff_A_iv4e9N5q4_0(.dout(w_dff_A_Vhb6DImv1_0),.din(w_dff_A_iv4e9N5q4_0),.clk(gclk));
	jdff dff_A_vjSqQ4gs1_0(.dout(w_Gid12_0[0]),.din(w_dff_A_vjSqQ4gs1_0),.clk(gclk));
	jdff dff_A_JuDPkQfu1_0(.dout(w_dff_A_vjSqQ4gs1_0),.din(w_dff_A_JuDPkQfu1_0),.clk(gclk));
	jdff dff_A_Qv375HHq5_0(.dout(w_dff_A_JuDPkQfu1_0),.din(w_dff_A_Qv375HHq5_0),.clk(gclk));
	jdff dff_A_QIqiZhg58_0(.dout(w_dff_A_Qv375HHq5_0),.din(w_dff_A_QIqiZhg58_0),.clk(gclk));
	jdff dff_A_BvHJu2zl3_0(.dout(w_dff_A_QIqiZhg58_0),.din(w_dff_A_BvHJu2zl3_0),.clk(gclk));
	jdff dff_A_Asr8THu82_0(.dout(w_dff_A_BvHJu2zl3_0),.din(w_dff_A_Asr8THu82_0),.clk(gclk));
	jdff dff_A_oOqD5JSR8_0(.dout(w_dff_A_Asr8THu82_0),.din(w_dff_A_oOqD5JSR8_0),.clk(gclk));
	jdff dff_A_6pNqEd4X3_0(.dout(w_dff_A_oOqD5JSR8_0),.din(w_dff_A_6pNqEd4X3_0),.clk(gclk));
	jdff dff_A_1YGnxI0q7_0(.dout(w_dff_A_6pNqEd4X3_0),.din(w_dff_A_1YGnxI0q7_0),.clk(gclk));
	jdff dff_B_R4HEtQGW7_1(.din(n90),.dout(w_dff_B_R4HEtQGW7_1),.clk(gclk));
	jdff dff_A_OTrU2NfY0_0(.dout(w_Gid7_0[0]),.din(w_dff_A_OTrU2NfY0_0),.clk(gclk));
	jdff dff_A_I9IxrMYY2_0(.dout(w_dff_A_OTrU2NfY0_0),.din(w_dff_A_I9IxrMYY2_0),.clk(gclk));
	jdff dff_A_4ojeLkYG9_0(.dout(w_dff_A_I9IxrMYY2_0),.din(w_dff_A_4ojeLkYG9_0),.clk(gclk));
	jdff dff_A_THSwPUtt4_0(.dout(w_dff_A_4ojeLkYG9_0),.din(w_dff_A_THSwPUtt4_0),.clk(gclk));
	jdff dff_A_n2MoqrZ97_0(.dout(w_dff_A_THSwPUtt4_0),.din(w_dff_A_n2MoqrZ97_0),.clk(gclk));
	jdff dff_A_l4Qsk1qB5_0(.dout(w_dff_A_n2MoqrZ97_0),.din(w_dff_A_l4Qsk1qB5_0),.clk(gclk));
	jdff dff_A_i4dMAA0L4_0(.dout(w_dff_A_l4Qsk1qB5_0),.din(w_dff_A_i4dMAA0L4_0),.clk(gclk));
	jdff dff_A_yMN71vaN3_0(.dout(w_dff_A_i4dMAA0L4_0),.din(w_dff_A_yMN71vaN3_0),.clk(gclk));
	jdff dff_A_DMwycXsd8_0(.dout(w_dff_A_yMN71vaN3_0),.din(w_dff_A_DMwycXsd8_0),.clk(gclk));
	jdff dff_A_94bBd39p7_0(.dout(w_Gid6_0[0]),.din(w_dff_A_94bBd39p7_0),.clk(gclk));
	jdff dff_A_hZhPAOVA3_0(.dout(w_dff_A_94bBd39p7_0),.din(w_dff_A_hZhPAOVA3_0),.clk(gclk));
	jdff dff_A_04XiGpaa8_0(.dout(w_dff_A_hZhPAOVA3_0),.din(w_dff_A_04XiGpaa8_0),.clk(gclk));
	jdff dff_A_AJHbVk5w4_0(.dout(w_dff_A_04XiGpaa8_0),.din(w_dff_A_AJHbVk5w4_0),.clk(gclk));
	jdff dff_A_hZcE0wOS9_0(.dout(w_dff_A_AJHbVk5w4_0),.din(w_dff_A_hZcE0wOS9_0),.clk(gclk));
	jdff dff_A_aOfOJiTD2_0(.dout(w_dff_A_hZcE0wOS9_0),.din(w_dff_A_aOfOJiTD2_0),.clk(gclk));
	jdff dff_A_OPBRgcvV5_0(.dout(w_dff_A_aOfOJiTD2_0),.din(w_dff_A_OPBRgcvV5_0),.clk(gclk));
	jdff dff_A_L0J8lgij4_0(.dout(w_dff_A_OPBRgcvV5_0),.din(w_dff_A_L0J8lgij4_0),.clk(gclk));
	jdff dff_A_7fxMyzXe9_0(.dout(w_dff_A_L0J8lgij4_0),.din(w_dff_A_7fxMyzXe9_0),.clk(gclk));
	jdff dff_A_caidO8Up4_0(.dout(w_Gid5_0[0]),.din(w_dff_A_caidO8Up4_0),.clk(gclk));
	jdff dff_A_YY7WWgQg2_0(.dout(w_dff_A_caidO8Up4_0),.din(w_dff_A_YY7WWgQg2_0),.clk(gclk));
	jdff dff_A_5FUYyccq4_0(.dout(w_dff_A_YY7WWgQg2_0),.din(w_dff_A_5FUYyccq4_0),.clk(gclk));
	jdff dff_A_CMouldip0_0(.dout(w_dff_A_5FUYyccq4_0),.din(w_dff_A_CMouldip0_0),.clk(gclk));
	jdff dff_A_XmXmT7pS5_0(.dout(w_dff_A_CMouldip0_0),.din(w_dff_A_XmXmT7pS5_0),.clk(gclk));
	jdff dff_A_LqB4KDHE2_0(.dout(w_dff_A_XmXmT7pS5_0),.din(w_dff_A_LqB4KDHE2_0),.clk(gclk));
	jdff dff_A_tngNbI3j8_0(.dout(w_dff_A_LqB4KDHE2_0),.din(w_dff_A_tngNbI3j8_0),.clk(gclk));
	jdff dff_A_JEOsdz1W0_0(.dout(w_dff_A_tngNbI3j8_0),.din(w_dff_A_JEOsdz1W0_0),.clk(gclk));
	jdff dff_A_f4JIbIaN0_0(.dout(w_dff_A_JEOsdz1W0_0),.din(w_dff_A_f4JIbIaN0_0),.clk(gclk));
	jdff dff_A_BhjqQ1Cs2_0(.dout(w_Gid4_0[0]),.din(w_dff_A_BhjqQ1Cs2_0),.clk(gclk));
	jdff dff_A_l71KpzS20_0(.dout(w_dff_A_BhjqQ1Cs2_0),.din(w_dff_A_l71KpzS20_0),.clk(gclk));
	jdff dff_A_VUtDisqQ5_0(.dout(w_dff_A_l71KpzS20_0),.din(w_dff_A_VUtDisqQ5_0),.clk(gclk));
	jdff dff_A_WaxHf69c0_0(.dout(w_dff_A_VUtDisqQ5_0),.din(w_dff_A_WaxHf69c0_0),.clk(gclk));
	jdff dff_A_OiVHDl0Z6_0(.dout(w_dff_A_WaxHf69c0_0),.din(w_dff_A_OiVHDl0Z6_0),.clk(gclk));
	jdff dff_A_Z7zZaQM37_0(.dout(w_dff_A_OiVHDl0Z6_0),.din(w_dff_A_Z7zZaQM37_0),.clk(gclk));
	jdff dff_A_HO71wEew0_0(.dout(w_dff_A_Z7zZaQM37_0),.din(w_dff_A_HO71wEew0_0),.clk(gclk));
	jdff dff_A_XRH2tvWv2_0(.dout(w_dff_A_HO71wEew0_0),.din(w_dff_A_XRH2tvWv2_0),.clk(gclk));
	jdff dff_A_D8w0sMRT0_0(.dout(w_dff_A_XRH2tvWv2_0),.din(w_dff_A_D8w0sMRT0_0),.clk(gclk));
endmodule

