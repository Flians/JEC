// Benchmark "c2670" written by ABC on Wed May 27 22:08:07 2020

module c2670 ( 
    G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
    G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
    G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
    G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
    G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
    G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
    G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119, G120,
    G123, G124, G125, G126, G127, G128, G129, G130, G131, G132, G135, G136,
    G137, G138, G139, G140, G141, G142, G169, G174, G177, G178, G179, G180,
    G181, G182, G183, G184, G185, G186, G189, G190, G191, G192, G193, G194,
    G195, G196, G197, G198, G199, G200, G201, G202, G203, G204, G205, G206,
    G207, G208, G209, G210, G211, G212, G213, G214, G215, G239, G240, G241,
    G242, G243, G244, G245, G246, G247, G248, G249, G250, G251, G252, G253,
    G254, G255, G256, G257, G262, G263, G264, G265, G266, G267, G268, G269,
    G270, G271, G272, G273, G274, G275, G276, G277, G278, G279, G452, G483,
    G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, G1384,
    G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, G2066,
    G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, G2106,
    G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20,
    G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36,
    G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56,
    G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74,
    G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90,
    G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105,
    G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
    G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132, G135,
    G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178, G179,
    G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192, G193,
    G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204, G205,
    G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239, G240,
    G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251, G252,
    G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267, G268,
    G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279, G452,
    G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348,
    G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996,
    G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105,
    G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474,
    G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire n381, n382, n383, n384, n385, n386, n388, n389, n390, n391, n394,
    n396, n398, n400, n401, n402, n403, n404, n405, n408, n409, n411, n412,
    n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
    n425, n426, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
    n438, n439, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
    n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
    n464, n465, n466, n467, n469, n470, n471, n472, n473, n474, n475, n476,
    n477, n479, n480, n481, n482, n483, n484, n487, n488, n489, n490, n491,
    n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n503, n504,
    n505, n506, n507, n509, n510, n512, n513, n514, n515, n516, n517, n518,
    n519, n520, n521, n525, n526, n527, n528, n529, n531, n532, n533, n534,
    n535, n536, n538, n539, n540, n541, n542, n543, n545, n546, n547, n548,
    n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n560, n561,
    n563, n565, n566, n567, n569, n570, n571, n572, n573, n574, n575, n576,
    n577, n578, n579, n580, n581, n583, n584, n585, n586, n587, n588, n589,
    n590, n591, n592, n593, n594, n595, n597, n598, n599, n600, n601, n602,
    n604, n605, n606, n607, n608, n609, n610, n611, n612, n614, n615, n616,
    n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
    n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
    n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
    n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
    n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
    n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
    n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
    n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
    n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
    n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
    n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
    n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
    n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
    n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
    n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
    n797, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
    n810, n811, n812, n813, n814, n815, n816, n818, n819, n820, n821, n822,
    n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n834, n835,
    n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
    n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
    n860, n861, n862, n863, n864, n865, n866, n867, n869, n870, n871, n872,
    n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n884, n885,
    n886, n887, n888, n889, n890, n891, n893, n894, n895, n896, n897, n898,
    n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
    n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
    n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
    n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
    n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
    n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
    n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
    n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
    n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
    n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
    n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
    n1026, n1027, n1028, n1029, n1032, n1033, n1034, n1035;
  jnot g000(.din(G44), .dout(G218));
  jnot g001(.din(G132), .dout(G219));
  jnot g002(.din(G82), .dout(G220));
  jnot g003(.din(G96), .dout(G221));
  jnot g004(.din(G69), .dout(G235));
  jnot g005(.din(G120), .dout(G236));
  jnot g006(.din(G57), .dout(G237));
  jnot g007(.din(G108), .dout(G238));
  jnot g008(.din(G2084), .dout(n381));
  jnot g009(.din(G2090), .dout(n382));
  jor  g010(.dina(n382), .dinb(n381), .dout(n383));
  jnot g011(.din(G2072), .dout(n384));
  jnot g012(.din(G2078), .dout(n385));
  jor  g013(.dina(n385), .dinb(n384), .dout(n386));
  jor  g014(.dina(n386), .dinb(n383), .dout(G158));
  jnot g015(.din(G15), .dout(n388));
  jnot g016(.din(G2), .dout(n389));
  jnot g017(.din(G661), .dout(n390));
  jor  g018(.dina(n390), .dinb(n389), .dout(n391));
  jor  g019(.dina(n391), .dinb(n388), .dout(G259));
  jand g020(.dina(G452), .dinb(G94), .dout(G173));
  jnot g021(.din(G7), .dout(n394));
  jor  g022(.dina(n390), .dinb(n394), .dout(G223));
  jnot g023(.din(G567), .dout(n396));
  jor  g024(.dina(G223), .dinb(n396), .dout(G234));
  jnot g025(.din(G2106), .dout(n398));
  jor  g026(.dina(G223), .dinb(n398), .dout(G217));
  jand g027(.dina(G108), .dinb(G69), .dout(n400));
  jand g028(.dina(G120), .dinb(G57), .dout(n401));
  jand g029(.dina(n401), .dinb(n400), .dout(n402));
  jand g030(.dina(G96), .dinb(G44), .dout(n403));
  jand g031(.dina(G132), .dinb(G82), .dout(n404));
  jand g032(.dina(n404), .dinb(n403), .dout(n405));
  jand g033(.dina(n405), .dinb(n402), .dout(G325));
  jnot g034(.din(G325), .dout(G261));
  jor  g035(.dina(n405), .dinb(n398), .dout(n408));
  jor  g036(.dina(n402), .dinb(n396), .dout(n409));
  jand g037(.dina(n409), .dinb(n408), .dout(G319));
  jnot g038(.din(G113), .dout(n411));
  jnot g039(.din(G2104), .dout(n412));
  jnot g040(.din(G2105), .dout(n413));
  jor  g041(.dina(n413), .dinb(n412), .dout(n414));
  jor  g042(.dina(n414), .dinb(n411), .dout(n415));
  jnot g043(.din(G101), .dout(n416));
  jor  g044(.dina(G2105), .dinb(n412), .dout(n417));
  jor  g045(.dina(n417), .dinb(n416), .dout(n418));
  jand g046(.dina(n418), .dinb(n415), .dout(n419));
  jnot g047(.din(G125), .dout(n420));
  jor  g048(.dina(n413), .dinb(G2104), .dout(n421));
  jor  g049(.dina(n421), .dinb(n420), .dout(n422));
  jnot g050(.din(G137), .dout(n423));
  jor  g051(.dina(G2105), .dinb(G2104), .dout(n424));
  jor  g052(.dina(n424), .dinb(n423), .dout(n425));
  jand g053(.dina(n425), .dinb(n422), .dout(n426));
  jand g054(.dina(n426), .dinb(n419), .dout(G160));
  jand g055(.dina(G2105), .dinb(G2104), .dout(n428));
  jand g056(.dina(n428), .dinb(G112), .dout(n429));
  jand g057(.dina(n413), .dinb(G2104), .dout(n430));
  jand g058(.dina(n430), .dinb(G100), .dout(n431));
  jor  g059(.dina(n431), .dinb(n429), .dout(n432));
  jnot g060(.din(n432), .dout(n433));
  jand g061(.dina(G2105), .dinb(n412), .dout(n434));
  jand g062(.dina(n434), .dinb(G124), .dout(n435));
  jnot g063(.din(n435), .dout(n436));
  jnot g064(.din(G136), .dout(n437));
  jor  g065(.dina(n424), .dinb(n437), .dout(n438));
  jand g066(.dina(n438), .dinb(n436), .dout(n439));
  jand g067(.dina(n439), .dinb(n433), .dout(G162));
  jnot g068(.din(G114), .dout(n441));
  jor  g069(.dina(n414), .dinb(n441), .dout(n442));
  jnot g070(.din(G102), .dout(n443));
  jor  g071(.dina(n417), .dinb(n443), .dout(n444));
  jand g072(.dina(n444), .dinb(n442), .dout(n445));
  jnot g073(.din(G126), .dout(n446));
  jor  g074(.dina(n421), .dinb(n446), .dout(n447));
  jnot g075(.din(G138), .dout(n448));
  jor  g076(.dina(n424), .dinb(n448), .dout(n449));
  jand g077(.dina(n449), .dinb(n447), .dout(n450));
  jand g078(.dina(n450), .dinb(n445), .dout(G164));
  jand g079(.dina(G651), .dinb(G543), .dout(n452));
  jand g080(.dina(n452), .dinb(G75), .dout(n453));
  jnot g081(.din(G651), .dout(n454));
  jand g082(.dina(n454), .dinb(G543), .dout(n455));
  jand g083(.dina(n455), .dinb(G50), .dout(n456));
  jor  g084(.dina(n456), .dinb(n453), .dout(n457));
  jnot g085(.din(n457), .dout(n458));
  jnot g086(.din(G543), .dout(n459));
  jand g087(.dina(G651), .dinb(n459), .dout(n460));
  jand g088(.dina(n460), .dinb(G62), .dout(n461));
  jnot g089(.din(n461), .dout(n462));
  jnot g090(.din(G88), .dout(n463));
  jand g091(.dina(n454), .dinb(n459), .dout(n464));
  jnot g092(.din(n464), .dout(n465));
  jor  g093(.dina(n465), .dinb(n463), .dout(n466));
  jand g094(.dina(n466), .dinb(n462), .dout(n467));
  jand g095(.dina(n467), .dinb(n458), .dout(G166));
  jand g096(.dina(n452), .dinb(G76), .dout(n469));
  jand g097(.dina(n455), .dinb(G51), .dout(n470));
  jor  g098(.dina(n470), .dinb(n469), .dout(n471));
  jnot g099(.din(n471), .dout(n472));
  jand g100(.dina(n460), .dinb(G63), .dout(n473));
  jnot g101(.din(n473), .dout(n474));
  jnot g102(.din(G89), .dout(n475));
  jor  g103(.dina(n465), .dinb(n475), .dout(n476));
  jand g104(.dina(n476), .dinb(n474), .dout(n477));
  jand g105(.dina(n477), .dinb(n472), .dout(G168));
  jand g106(.dina(n452), .dinb(G77), .dout(n479));
  jand g107(.dina(n455), .dinb(G52), .dout(n480));
  jor  g108(.dina(n480), .dinb(n479), .dout(n481));
  jand g109(.dina(n460), .dinb(G64), .dout(n482));
  jand g110(.dina(n464), .dinb(G90), .dout(n483));
  jor  g111(.dina(n483), .dinb(n482), .dout(n484));
  jor  g112(.dina(n484), .dinb(n481), .dout(G301));
  jnot g113(.din(G301), .dout(G171));
  jnot g114(.din(G860), .dout(n487));
  jand g115(.dina(n452), .dinb(G68), .dout(n488));
  jnot g116(.din(n488), .dout(n489));
  jnot g117(.din(G43), .dout(n490));
  jnot g118(.din(n455), .dout(n491));
  jor  g119(.dina(n491), .dinb(n490), .dout(n492));
  jand g120(.dina(n492), .dinb(n489), .dout(n493));
  jnot g121(.din(G56), .dout(n494));
  jnot g122(.din(n460), .dout(n495));
  jor  g123(.dina(n495), .dinb(n494), .dout(n496));
  jnot g124(.din(G81), .dout(n497));
  jor  g125(.dina(n465), .dinb(n497), .dout(n498));
  jand g126(.dina(n498), .dinb(n496), .dout(n499));
  jand g127(.dina(n499), .dinb(n493), .dout(n500));
  jnot g128(.din(n500), .dout(n501));
  jor  g129(.dina(n501), .dinb(n487), .dout(G153));
  jnot g130(.din(G319), .dout(n503));
  jnot g131(.din(G36), .dout(n504));
  jnot g132(.din(G483), .dout(n505));
  jor  g133(.dina(n390), .dinb(n505), .dout(n506));
  jor  g134(.dina(n506), .dinb(n504), .dout(n507));
  jor  g135(.dina(n507), .dinb(n503), .dout(G176));
  jand g136(.dina(G3), .dinb(G1), .dout(n509));
  jor  g137(.dina(n509), .dinb(n506), .dout(n510));
  jor  g138(.dina(n510), .dinb(n503), .dout(G188));
  jand g139(.dina(n452), .dinb(G78), .dout(n512));
  jand g140(.dina(n455), .dinb(G53), .dout(n513));
  jor  g141(.dina(n513), .dinb(n512), .dout(n514));
  jnot g142(.din(n514), .dout(n515));
  jand g143(.dina(n460), .dinb(G65), .dout(n516));
  jnot g144(.din(n516), .dout(n517));
  jnot g145(.din(G91), .dout(n518));
  jor  g146(.dina(n465), .dinb(n518), .dout(n519));
  jand g147(.dina(n519), .dinb(n517), .dout(n520));
  jand g148(.dina(n520), .dinb(n515), .dout(n521));
  jnot g149(.din(n521), .dout(G299));
  jnot g150(.din(G168), .dout(G286));
  jnot g151(.din(G166), .dout(G303));
  jand g152(.dina(n464), .dinb(G87), .dout(n525));
  jor  g153(.dina(n525), .dinb(n460), .dout(n526));
  jand g154(.dina(n455), .dinb(G49), .dout(n527));
  jand g155(.dina(n452), .dinb(G74), .dout(n528));
  jor  g156(.dina(n528), .dinb(n527), .dout(n529));
  jor  g157(.dina(n529), .dinb(n526), .dout(G288));
  jand g158(.dina(n452), .dinb(G73), .dout(n531));
  jand g159(.dina(n455), .dinb(G48), .dout(n532));
  jor  g160(.dina(n532), .dinb(n531), .dout(n533));
  jand g161(.dina(n460), .dinb(G61), .dout(n534));
  jand g162(.dina(n464), .dinb(G86), .dout(n535));
  jor  g163(.dina(n535), .dinb(n534), .dout(n536));
  jor  g164(.dina(n536), .dinb(n533), .dout(G305));
  jand g165(.dina(n452), .dinb(G72), .dout(n538));
  jand g166(.dina(n455), .dinb(G47), .dout(n539));
  jor  g167(.dina(n539), .dinb(n538), .dout(n540));
  jand g168(.dina(n460), .dinb(G60), .dout(n541));
  jand g169(.dina(n464), .dinb(G85), .dout(n542));
  jor  g170(.dina(n542), .dinb(n541), .dout(n543));
  jor  g171(.dina(n543), .dinb(n540), .dout(G290));
  jnot g172(.din(G868), .dout(n545));
  jand g173(.dina(n452), .dinb(G79), .dout(n546));
  jand g174(.dina(n455), .dinb(G54), .dout(n547));
  jor  g175(.dina(n547), .dinb(n546), .dout(n548));
  jnot g176(.din(n548), .dout(n549));
  jand g177(.dina(n460), .dinb(G66), .dout(n550));
  jnot g178(.din(n550), .dout(n551));
  jnot g179(.din(G92), .dout(n552));
  jor  g180(.dina(n465), .dinb(n552), .dout(n553));
  jand g181(.dina(n553), .dinb(n551), .dout(n554));
  jand g182(.dina(n554), .dinb(n549), .dout(n555));
  jnot g183(.din(n555), .dout(n556));
  jand g184(.dina(n556), .dinb(n545), .dout(n557));
  jand g185(.dina(G301), .dinb(G868), .dout(n558));
  jor  g186(.dina(n558), .dinb(n557), .dout(G284));
  jand g187(.dina(G299), .dinb(n545), .dout(n560));
  jand g188(.dina(G286), .dinb(G868), .dout(n561));
  jor  g189(.dina(n561), .dinb(n560), .dout(G297));
  jand g190(.dina(n487), .dinb(G559), .dout(n563));
  jor  g191(.dina(n563), .dinb(n556), .dout(G148));
  jor  g192(.dina(n556), .dinb(G559), .dout(n565));
  jand g193(.dina(n565), .dinb(G868), .dout(n566));
  jand g194(.dina(n501), .dinb(n545), .dout(n567));
  jor  g195(.dina(n567), .dinb(n566), .dout(G282));
  jand g196(.dina(n428), .dinb(G111), .dout(n569));
  jand g197(.dina(n430), .dinb(G99), .dout(n570));
  jor  g198(.dina(n570), .dinb(n569), .dout(n571));
  jand g199(.dina(n434), .dinb(G123), .dout(n572));
  jand g200(.dina(n413), .dinb(n412), .dout(n573));
  jand g201(.dina(n573), .dinb(G135), .dout(n574));
  jor  g202(.dina(n574), .dinb(n572), .dout(n575));
  jor  g203(.dina(n575), .dinb(n571), .dout(n576));
  jand g204(.dina(n576), .dinb(G2096), .dout(n577));
  jnot g205(.din(G2096), .dout(n578));
  jnot g206(.din(n576), .dout(n579));
  jand g207(.dina(n579), .dinb(n578), .dout(n580));
  jor  g208(.dina(n580), .dinb(G2100), .dout(n581));
  jor  g209(.dina(n581), .dinb(n577), .dout(G156));
  jxor g210(.dina(G2446), .dinb(G2443), .dout(n583));
  jnot g211(.din(n583), .dout(n584));
  jxor g212(.dina(G2454), .dinb(G2451), .dout(n585));
  jxor g213(.dina(G1348), .dinb(G1341), .dout(n586));
  jxor g214(.dina(n586), .dinb(n585), .dout(n587));
  jxor g215(.dina(G2430), .dinb(G2427), .dout(n588));
  jxor g216(.dina(G2438), .dinb(G2435), .dout(n589));
  jxor g217(.dina(n589), .dinb(n588), .dout(n590));
  jxor g218(.dina(n590), .dinb(n587), .dout(n591));
  jand g219(.dina(n591), .dinb(n584), .dout(n592));
  jnot g220(.din(n592), .dout(n593));
  jor  g221(.dina(n591), .dinb(n584), .dout(n594));
  jand g222(.dina(n594), .dinb(G14), .dout(n595));
  jand g223(.dina(n595), .dinb(n593), .dout(G401));
  jxor g224(.dina(G2100), .dinb(n578), .dout(n597));
  jxor g225(.dina(G2078), .dinb(G2072), .dout(n598));
  jxor g226(.dina(G2090), .dinb(G2084), .dout(n599));
  jxor g227(.dina(G2678), .dinb(G2067), .dout(n600));
  jxor g228(.dina(n600), .dinb(n599), .dout(n601));
  jxor g229(.dina(n601), .dinb(n598), .dout(n602));
  jxor g230(.dina(n602), .dinb(n597), .dout(G227));
  jxor g231(.dina(G1986), .dinb(G1981), .dout(n604));
  jxor g232(.dina(G1966), .dinb(G1961), .dout(n605));
  jxor g233(.dina(n605), .dinb(n604), .dout(n606));
  jxor g234(.dina(G2474), .dinb(G1956), .dout(n607));
  jxor g235(.dina(G1976), .dinb(G1971), .dout(n608));
  jxor g236(.dina(n608), .dinb(n607), .dout(n609));
  jnot g237(.din(G1991), .dout(n610));
  jxor g238(.dina(G1996), .dinb(n610), .dout(n611));
  jxor g239(.dina(n611), .dinb(n609), .dout(n612));
  jxor g240(.dina(n612), .dinb(n606), .dout(G229));
  jand g241(.dina(G290), .dinb(G16), .dout(n614));
  jnot g242(.din(G16), .dout(n615));
  jand g243(.dina(G24), .dinb(n615), .dout(n616));
  jor  g244(.dina(n616), .dinb(n614), .dout(n617));
  jand g245(.dina(n617), .dinb(G1986), .dout(n618));
  jnot g246(.din(n618), .dout(n619));
  jor  g247(.dina(G34), .dinb(G29), .dout(n620));
  jnot g248(.din(n620), .dout(n621));
  jand g249(.dina(G160), .dinb(G29), .dout(n622));
  jor  g250(.dina(n622), .dinb(n621), .dout(n623));
  jand g251(.dina(n623), .dinb(n381), .dout(n624));
  jnot g252(.din(n624), .dout(n625));
  jor  g253(.dina(n617), .dinb(G1986), .dout(n626));
  jand g254(.dina(n626), .dinb(n625), .dout(n627));
  jand g255(.dina(n627), .dinb(n619), .dout(n628));
  jor  g256(.dina(n623), .dinb(n381), .dout(n629));
  jor  g257(.dina(G32), .dinb(G29), .dout(n630));
  jand g258(.dina(n428), .dinb(G117), .dout(n631));
  jand g259(.dina(n430), .dinb(G105), .dout(n632));
  jor  g260(.dina(n632), .dinb(n631), .dout(n633));
  jnot g261(.din(n633), .dout(n634));
  jand g262(.dina(n434), .dinb(G129), .dout(n635));
  jnot g263(.din(n635), .dout(n636));
  jnot g264(.din(G141), .dout(n637));
  jor  g265(.dina(n424), .dinb(n637), .dout(n638));
  jand g266(.dina(n638), .dinb(n636), .dout(n639));
  jand g267(.dina(n639), .dinb(n634), .dout(n640));
  jand g268(.dina(n640), .dinb(G29), .dout(n641));
  jnot g269(.din(n641), .dout(n642));
  jand g270(.dina(n642), .dinb(n630), .dout(n643));
  jand g271(.dina(n643), .dinb(G1996), .dout(n644));
  jnot g272(.din(n644), .dout(n645));
  jand g273(.dina(n645), .dinb(n629), .dout(n646));
  jnot g274(.din(G1966), .dout(n647));
  jor  g275(.dina(G21), .dinb(G16), .dout(n648));
  jand g276(.dina(G168), .dinb(G16), .dout(n649));
  jnot g277(.din(n649), .dout(n650));
  jand g278(.dina(n650), .dinb(n648), .dout(n651));
  jnot g279(.din(n651), .dout(n652));
  jand g280(.dina(n652), .dinb(n647), .dout(n653));
  jor  g281(.dina(G29), .dinb(G27), .dout(n654));
  jnot g282(.din(n654), .dout(n655));
  jand g283(.dina(G164), .dinb(G29), .dout(n656));
  jor  g284(.dina(n656), .dinb(n655), .dout(n657));
  jand g285(.dina(n657), .dinb(n385), .dout(n658));
  jor  g286(.dina(n658), .dinb(n653), .dout(n659));
  jnot g287(.din(n659), .dout(n660));
  jand g288(.dina(n660), .dinb(n646), .dout(n661));
  jor  g289(.dina(G35), .dinb(G29), .dout(n662));
  jand g290(.dina(G162), .dinb(G29), .dout(n663));
  jnot g291(.din(n663), .dout(n664));
  jand g292(.dina(n664), .dinb(n662), .dout(n665));
  jnot g293(.din(n665), .dout(n666));
  jand g294(.dina(n666), .dinb(n382), .dout(n667));
  jor  g295(.dina(G29), .dinb(G26), .dout(n668));
  jand g296(.dina(n428), .dinb(G116), .dout(n669));
  jand g297(.dina(n430), .dinb(G104), .dout(n670));
  jor  g298(.dina(n670), .dinb(n669), .dout(n671));
  jnot g299(.din(n671), .dout(n672));
  jand g300(.dina(n434), .dinb(G128), .dout(n673));
  jnot g301(.din(n673), .dout(n674));
  jnot g302(.din(G140), .dout(n675));
  jor  g303(.dina(n424), .dinb(n675), .dout(n676));
  jand g304(.dina(n676), .dinb(n674), .dout(n677));
  jand g305(.dina(n677), .dinb(n672), .dout(n678));
  jand g306(.dina(n678), .dinb(G29), .dout(n679));
  jnot g307(.din(n679), .dout(n680));
  jand g308(.dina(n680), .dinb(n668), .dout(n681));
  jand g309(.dina(n681), .dinb(G2067), .dout(n682));
  jor  g310(.dina(n682), .dinb(n667), .dout(n683));
  jnot g311(.din(G1348), .dout(n684));
  jor  g312(.dina(G16), .dinb(G4), .dout(n685));
  jand g313(.dina(n555), .dinb(G16), .dout(n686));
  jnot g314(.din(n686), .dout(n687));
  jand g315(.dina(n687), .dinb(n685), .dout(n688));
  jnot g316(.din(n688), .dout(n689));
  jand g317(.dina(n689), .dinb(n684), .dout(n690));
  jnot g318(.din(G1981), .dout(n691));
  jand g319(.dina(G305), .dinb(G16), .dout(n692));
  jand g320(.dina(n615), .dinb(G6), .dout(n693));
  jor  g321(.dina(n693), .dinb(n692), .dout(n694));
  jnot g322(.din(n694), .dout(n695));
  jand g323(.dina(n695), .dinb(n691), .dout(n696));
  jor  g324(.dina(n696), .dinb(n690), .dout(n697));
  jor  g325(.dina(n697), .dinb(n683), .dout(n698));
  jnot g326(.din(n698), .dout(n699));
  jand g327(.dina(n699), .dinb(n661), .dout(n700));
  jand g328(.dina(n700), .dinb(n628), .dout(n701));
  jor  g329(.dina(G171), .dinb(n615), .dout(n702));
  jnot g330(.din(G5), .dout(n703));
  jor  g331(.dina(G16), .dinb(n703), .dout(n704));
  jand g332(.dina(n704), .dinb(n702), .dout(n705));
  jxor g333(.dina(n705), .dinb(G1961), .dout(n706));
  jnot g334(.din(n706), .dout(n707));
  jor  g335(.dina(G29), .dinb(G25), .dout(n708));
  jnot g336(.din(G29), .dout(n709));
  jand g337(.dina(n428), .dinb(G107), .dout(n710));
  jand g338(.dina(n430), .dinb(G95), .dout(n711));
  jor  g339(.dina(n711), .dinb(n710), .dout(n712));
  jand g340(.dina(n434), .dinb(G119), .dout(n713));
  jand g341(.dina(n573), .dinb(G131), .dout(n714));
  jor  g342(.dina(n714), .dinb(n713), .dout(n715));
  jor  g343(.dina(n715), .dinb(n712), .dout(n716));
  jor  g344(.dina(n716), .dinb(n709), .dout(n717));
  jand g345(.dina(n717), .dinb(n708), .dout(n718));
  jxor g346(.dina(n718), .dinb(n610), .dout(n719));
  jnot g347(.din(n719), .dout(n720));
  jor  g348(.dina(n657), .dinb(n385), .dout(n721));
  jand g349(.dina(n579), .dinb(G29), .dout(n722));
  jor  g350(.dina(G29), .dinb(G28), .dout(n723));
  jand g351(.dina(n723), .dinb(G11), .dout(n724));
  jnot g352(.din(n724), .dout(n725));
  jor  g353(.dina(n725), .dinb(n722), .dout(n726));
  jnot g354(.din(n726), .dout(n727));
  jand g355(.dina(n727), .dinb(n721), .dout(n728));
  jand g356(.dina(n728), .dinb(n720), .dout(n729));
  jand g357(.dina(n729), .dinb(n707), .dout(n730));
  jor  g358(.dina(G33), .dinb(G29), .dout(n731));
  jand g359(.dina(n428), .dinb(G115), .dout(n732));
  jand g360(.dina(n430), .dinb(G103), .dout(n733));
  jor  g361(.dina(n733), .dinb(n732), .dout(n734));
  jnot g362(.din(n734), .dout(n735));
  jand g363(.dina(n434), .dinb(G127), .dout(n736));
  jnot g364(.din(n736), .dout(n737));
  jnot g365(.din(G139), .dout(n738));
  jor  g366(.dina(n424), .dinb(n738), .dout(n739));
  jand g367(.dina(n739), .dinb(n737), .dout(n740));
  jand g368(.dina(n740), .dinb(n735), .dout(n741));
  jand g369(.dina(n741), .dinb(G29), .dout(n742));
  jnot g370(.din(n742), .dout(n743));
  jand g371(.dina(n743), .dinb(n731), .dout(n744));
  jor  g372(.dina(n744), .dinb(G2072), .dout(n745));
  jor  g373(.dina(G20), .dinb(G16), .dout(n746));
  jand g374(.dina(n521), .dinb(G16), .dout(n747));
  jnot g375(.din(n747), .dout(n748));
  jand g376(.dina(n748), .dinb(n746), .dout(n749));
  jor  g377(.dina(n749), .dinb(G1956), .dout(n750));
  jand g378(.dina(n750), .dinb(n745), .dout(n751));
  jor  g379(.dina(G22), .dinb(G16), .dout(n752));
  jand g380(.dina(G166), .dinb(G16), .dout(n753));
  jnot g381(.din(n753), .dout(n754));
  jand g382(.dina(n754), .dinb(n752), .dout(n755));
  jor  g383(.dina(n755), .dinb(G1971), .dout(n756));
  jand g384(.dina(n665), .dinb(G2090), .dout(n757));
  jnot g385(.din(n757), .dout(n758));
  jand g386(.dina(n758), .dinb(n756), .dout(n759));
  jand g387(.dina(n759), .dinb(n751), .dout(n760));
  jor  g388(.dina(n681), .dinb(G2067), .dout(n761));
  jand g389(.dina(n694), .dinb(G1981), .dout(n762));
  jnot g390(.din(n762), .dout(n763));
  jand g391(.dina(n763), .dinb(n761), .dout(n764));
  jand g392(.dina(n651), .dinb(G1966), .dout(n765));
  jand g393(.dina(n755), .dinb(G1971), .dout(n766));
  jor  g394(.dina(n766), .dinb(n765), .dout(n767));
  jnot g395(.din(n767), .dout(n768));
  jand g396(.dina(n768), .dinb(n764), .dout(n769));
  jand g397(.dina(n769), .dinb(n760), .dout(n770));
  jnot g398(.din(G1976), .dout(n771));
  jand g399(.dina(G288), .dinb(G16), .dout(n772));
  jand g400(.dina(G23), .dinb(n615), .dout(n773));
  jor  g401(.dina(n773), .dinb(n772), .dout(n774));
  jnot g402(.din(n774), .dout(n775));
  jand g403(.dina(n775), .dinb(n771), .dout(n776));
  jnot g404(.din(n776), .dout(n777));
  jor  g405(.dina(n643), .dinb(G1996), .dout(n778));
  jand g406(.dina(n778), .dinb(n777), .dout(n779));
  jand g407(.dina(n749), .dinb(G1956), .dout(n780));
  jand g408(.dina(n774), .dinb(G1976), .dout(n781));
  jor  g409(.dina(n781), .dinb(n780), .dout(n782));
  jnot g410(.din(n782), .dout(n783));
  jand g411(.dina(n783), .dinb(n779), .dout(n784));
  jor  g412(.dina(G19), .dinb(G16), .dout(n785));
  jor  g413(.dina(n501), .dinb(n615), .dout(n786));
  jand g414(.dina(n786), .dinb(n785), .dout(n787));
  jxor g415(.dina(n787), .dinb(G1341), .dout(n788));
  jnot g416(.din(n788), .dout(n789));
  jand g417(.dina(n688), .dinb(G1348), .dout(n790));
  jand g418(.dina(n744), .dinb(G2072), .dout(n791));
  jor  g419(.dina(n791), .dinb(n790), .dout(n792));
  jor  g420(.dina(n792), .dinb(n789), .dout(n793));
  jnot g421(.din(n793), .dout(n794));
  jand g422(.dina(n794), .dinb(n784), .dout(n795));
  jand g423(.dina(n795), .dinb(n770), .dout(n796));
  jand g424(.dina(n796), .dinb(n730), .dout(n797));
  jand g425(.dina(n797), .dinb(n701), .dout(G311));
  jnot g426(.din(n628), .dout(n799));
  jnot g427(.din(n646), .dout(n800));
  jor  g428(.dina(n659), .dinb(n800), .dout(n801));
  jor  g429(.dina(n698), .dinb(n801), .dout(n802));
  jor  g430(.dina(n802), .dinb(n799), .dout(n803));
  jnot g431(.din(n730), .dout(n804));
  jnot g432(.din(n751), .dout(n805));
  jnot g433(.din(n756), .dout(n806));
  jor  g434(.dina(n757), .dinb(n806), .dout(n807));
  jor  g435(.dina(n807), .dinb(n805), .dout(n808));
  jnot g436(.din(n764), .dout(n809));
  jor  g437(.dina(n767), .dinb(n809), .dout(n810));
  jor  g438(.dina(n810), .dinb(n808), .dout(n811));
  jnot g439(.din(n779), .dout(n812));
  jor  g440(.dina(n782), .dinb(n812), .dout(n813));
  jor  g441(.dina(n793), .dinb(n813), .dout(n814));
  jor  g442(.dina(n814), .dinb(n811), .dout(n815));
  jor  g443(.dina(n815), .dinb(n804), .dout(n816));
  jor  g444(.dina(n816), .dinb(n803), .dout(G150));
  jnot g445(.din(n563), .dout(n818));
  jor  g446(.dina(n818), .dinb(n556), .dout(n819));
  jand g447(.dina(n819), .dinb(G153), .dout(n820));
  jand g448(.dina(n452), .dinb(G80), .dout(n821));
  jnot g449(.din(n821), .dout(n822));
  jnot g450(.din(G55), .dout(n823));
  jor  g451(.dina(n491), .dinb(n823), .dout(n824));
  jand g452(.dina(n824), .dinb(n822), .dout(n825));
  jnot g453(.din(G67), .dout(n826));
  jor  g454(.dina(n495), .dinb(n826), .dout(n827));
  jnot g455(.din(G93), .dout(n828));
  jor  g456(.dina(n465), .dinb(n828), .dout(n829));
  jand g457(.dina(n829), .dinb(n827), .dout(n830));
  jand g458(.dina(n830), .dinb(n825), .dout(n831));
  jxor g459(.dina(n831), .dinb(n500), .dout(n832));
  jxor g460(.dina(n832), .dinb(n820), .dout(G145));
  jand g461(.dina(n428), .dinb(G113), .dout(n834));
  jand g462(.dina(n430), .dinb(G101), .dout(n835));
  jor  g463(.dina(n835), .dinb(n834), .dout(n836));
  jand g464(.dina(n434), .dinb(G125), .dout(n837));
  jand g465(.dina(n573), .dinb(G137), .dout(n838));
  jor  g466(.dina(n838), .dinb(n837), .dout(n839));
  jor  g467(.dina(n839), .dinb(n836), .dout(n840));
  jxor g468(.dina(G162), .dinb(n840), .dout(n841));
  jxor g469(.dina(n841), .dinb(n579), .dout(n842));
  jxor g470(.dina(n716), .dinb(n678), .dout(n843));
  jand g471(.dina(n428), .dinb(G118), .dout(n844));
  jand g472(.dina(n430), .dinb(G106), .dout(n845));
  jor  g473(.dina(n845), .dinb(n844), .dout(n846));
  jand g474(.dina(n434), .dinb(G130), .dout(n847));
  jand g475(.dina(n573), .dinb(G142), .dout(n848));
  jor  g476(.dina(n848), .dinb(n847), .dout(n849));
  jor  g477(.dina(n849), .dinb(n846), .dout(n850));
  jand g478(.dina(n428), .dinb(G114), .dout(n851));
  jand g479(.dina(n430), .dinb(G102), .dout(n852));
  jor  g480(.dina(n852), .dinb(n851), .dout(n853));
  jand g481(.dina(n434), .dinb(G126), .dout(n854));
  jand g482(.dina(n573), .dinb(G138), .dout(n855));
  jor  g483(.dina(n855), .dinb(n854), .dout(n856));
  jor  g484(.dina(n856), .dinb(n853), .dout(n857));
  jxor g485(.dina(n640), .dinb(n857), .dout(n858));
  jxor g486(.dina(n858), .dinb(n741), .dout(n859));
  jxor g487(.dina(n859), .dinb(n850), .dout(n860));
  jxor g488(.dina(n860), .dinb(n843), .dout(n861));
  jnot g489(.din(n861), .dout(n862));
  jand g490(.dina(n862), .dinb(n842), .dout(n863));
  jnot g491(.din(n842), .dout(n864));
  jand g492(.dina(n861), .dinb(n864), .dout(n865));
  jor  g493(.dina(n865), .dinb(G37), .dout(n866));
  jor  g494(.dina(n866), .dinb(n863), .dout(n867));
  jnot g495(.din(n867), .dout(G395));
  jxor g496(.dina(G305), .dinb(G166), .dout(n869));
  jnot g497(.din(G288), .dout(n870));
  jxor g498(.dina(G290), .dinb(n870), .dout(n871));
  jxor g499(.dina(n871), .dinb(n869), .dout(n872));
  jxor g500(.dina(n832), .dinb(G299), .dout(n873));
  jor  g501(.dina(n873), .dinb(n565), .dout(n874));
  jnot g502(.din(n565), .dout(n875));
  jxor g503(.dina(n873), .dinb(n555), .dout(n876));
  jor  g504(.dina(n876), .dinb(n875), .dout(n877));
  jand g505(.dina(n877), .dinb(n874), .dout(n878));
  jxor g506(.dina(n878), .dinb(n872), .dout(n879));
  jand g507(.dina(n879), .dinb(G868), .dout(n880));
  jnot g508(.din(n831), .dout(n881));
  jand g509(.dina(n881), .dinb(n545), .dout(n882));
  jor  g510(.dina(n882), .dinb(n880), .dout(G295));
  jnot g511(.din(n872), .dout(n884));
  jxor g512(.dina(G301), .dinb(G168), .dout(n885));
  jxor g513(.dina(n885), .dinb(n876), .dout(n886));
  jand g514(.dina(n886), .dinb(n884), .dout(n887));
  jnot g515(.din(n887), .dout(n888));
  jnot g516(.din(G37), .dout(n889));
  jor  g517(.dina(n886), .dinb(n884), .dout(n890));
  jand g518(.dina(n890), .dinb(n889), .dout(n891));
  jand g519(.dina(n891), .dinb(n888), .dout(G397));
  jnot g520(.din(G1341), .dout(n893));
  jnot g521(.din(G1384), .dout(n894));
  jand g522(.dina(n857), .dinb(n894), .dout(n895));
  jand g523(.dina(G160), .dinb(G40), .dout(n896));
  jand g524(.dina(n896), .dinb(n895), .dout(n897));
  jor  g525(.dina(n897), .dinb(n893), .dout(n898));
  jnot g526(.din(G1996), .dout(n899));
  jor  g527(.dina(G164), .dinb(G1384), .dout(n900));
  jnot g528(.din(G40), .dout(n901));
  jor  g529(.dina(n840), .dinb(n901), .dout(n902));
  jor  g530(.dina(n902), .dinb(n900), .dout(n903));
  jor  g531(.dina(n903), .dinb(n899), .dout(n904));
  jand g532(.dina(n904), .dinb(n500), .dout(n905));
  jand g533(.dina(n905), .dinb(n898), .dout(n906));
  jor  g534(.dina(n906), .dinb(n555), .dout(n907));
  jor  g535(.dina(n897), .dinb(n684), .dout(n908));
  jnot g536(.din(G2067), .dout(n909));
  jor  g537(.dina(n903), .dinb(n909), .dout(n910));
  jand g538(.dina(n910), .dinb(n908), .dout(n911));
  jand g539(.dina(n911), .dinb(n907), .dout(n912));
  jnot g540(.din(G1956), .dout(n913));
  jor  g541(.dina(n897), .dinb(n913), .dout(n914));
  jor  g542(.dina(n903), .dinb(n384), .dout(n915));
  jand g543(.dina(n915), .dinb(n914), .dout(n916));
  jand g544(.dina(n916), .dinb(n521), .dout(n917));
  jand g545(.dina(n906), .dinb(n555), .dout(n918));
  jor  g546(.dina(n918), .dinb(n917), .dout(n919));
  jor  g547(.dina(n919), .dinb(n912), .dout(n920));
  jnot g548(.din(G1971), .dout(n921));
  jor  g549(.dina(n897), .dinb(n921), .dout(n922));
  jor  g550(.dina(n903), .dinb(n382), .dout(n923));
  jand g551(.dina(n923), .dinb(G8), .dout(n924));
  jand g552(.dina(n924), .dinb(n922), .dout(n925));
  jnot g553(.din(G8), .dout(n926));
  jor  g554(.dina(G166), .dinb(n926), .dout(n927));
  jor  g555(.dina(n927), .dinb(n925), .dout(n928));
  jand g556(.dina(n903), .dinb(G1971), .dout(n929));
  jand g557(.dina(n897), .dinb(G2090), .dout(n930));
  jor  g558(.dina(n930), .dinb(n926), .dout(n931));
  jor  g559(.dina(n931), .dinb(n929), .dout(n932));
  jor  g560(.dina(n932), .dinb(G303), .dout(n933));
  jand g561(.dina(n933), .dinb(n928), .dout(n934));
  jand g562(.dina(n691), .dinb(G8), .dout(n935));
  jnot g563(.din(n935), .dout(n936));
  jor  g564(.dina(n936), .dinb(G305), .dout(n937));
  jor  g565(.dina(n937), .dinb(n897), .dout(n938));
  jnot g566(.din(G305), .dout(n939));
  jor  g567(.dina(n691), .dinb(n926), .dout(n940));
  jor  g568(.dina(n940), .dinb(n939), .dout(n941));
  jor  g569(.dina(n941), .dinb(n897), .dout(n942));
  jand g570(.dina(n942), .dinb(n938), .dout(n943));
  jand g571(.dina(n771), .dinb(G8), .dout(n944));
  jnot g572(.din(n944), .dout(n945));
  jor  g573(.dina(n945), .dinb(G288), .dout(n946));
  jor  g574(.dina(n946), .dinb(n897), .dout(n947));
  jor  g575(.dina(n771), .dinb(n926), .dout(n948));
  jor  g576(.dina(n948), .dinb(n870), .dout(n949));
  jor  g577(.dina(n949), .dinb(n897), .dout(n950));
  jand g578(.dina(n950), .dinb(n947), .dout(n951));
  jand g579(.dina(n951), .dinb(n943), .dout(n952));
  jand g580(.dina(n952), .dinb(n934), .dout(n953));
  jor  g581(.dina(n897), .dinb(n647), .dout(n954));
  jor  g582(.dina(n903), .dinb(n381), .dout(n955));
  jand g583(.dina(n955), .dinb(G8), .dout(n956));
  jand g584(.dina(n956), .dinb(n954), .dout(n957));
  jor  g585(.dina(G168), .dinb(n926), .dout(n958));
  jor  g586(.dina(n958), .dinb(n957), .dout(n959));
  jand g587(.dina(n903), .dinb(G1966), .dout(n960));
  jand g588(.dina(n897), .dinb(G2084), .dout(n961));
  jor  g589(.dina(n961), .dinb(n926), .dout(n962));
  jor  g590(.dina(n962), .dinb(n960), .dout(n963));
  jor  g591(.dina(n963), .dinb(G286), .dout(n964));
  jand g592(.dina(n964), .dinb(n959), .dout(n965));
  jnot g593(.din(G1961), .dout(n966));
  jor  g594(.dina(n897), .dinb(n966), .dout(n967));
  jor  g595(.dina(n903), .dinb(n385), .dout(n968));
  jand g596(.dina(n968), .dinb(n967), .dout(n969));
  jor  g597(.dina(n969), .dinb(G171), .dout(n970));
  jand g598(.dina(n903), .dinb(G1961), .dout(n971));
  jand g599(.dina(n897), .dinb(G2078), .dout(n972));
  jor  g600(.dina(n972), .dinb(n971), .dout(n973));
  jor  g601(.dina(n973), .dinb(G301), .dout(n974));
  jor  g602(.dina(n916), .dinb(n521), .dout(n975));
  jand g603(.dina(n975), .dinb(n974), .dout(n976));
  jand g604(.dina(n976), .dinb(n970), .dout(n977));
  jand g605(.dina(n977), .dinb(n965), .dout(n978));
  jand g606(.dina(n978), .dinb(n953), .dout(n979));
  jand g607(.dina(n979), .dinb(n920), .dout(n980));
  jnot g608(.din(n974), .dout(n981));
  jand g609(.dina(n981), .dinb(n965), .dout(n982));
  jand g610(.dina(n982), .dinb(n953), .dout(n983));
  jand g611(.dina(n957), .dinb(G168), .dout(n984));
  jand g612(.dina(n984), .dinb(n952), .dout(n985));
  jand g613(.dina(n985), .dinb(n934), .dout(n986));
  jand g614(.dina(n925), .dinb(G166), .dout(n987));
  jand g615(.dina(n952), .dinb(n987), .dout(n988));
  jnot g616(.din(n938), .dout(n989));
  jnot g617(.din(n947), .dout(n990));
  jand g618(.dina(n990), .dinb(n942), .dout(n991));
  jor  g619(.dina(n991), .dinb(n989), .dout(n992));
  jor  g620(.dina(n992), .dinb(n988), .dout(n993));
  jor  g621(.dina(n993), .dinb(n986), .dout(n994));
  jor  g622(.dina(n994), .dinb(n983), .dout(n995));
  jor  g623(.dina(n995), .dinb(n980), .dout(n996));
  jand g624(.dina(n896), .dinb(n900), .dout(n997));
  jand g625(.dina(n678), .dinb(n909), .dout(n998));
  jand g626(.dina(n998), .dinb(n997), .dout(n999));
  jnot g627(.din(n999), .dout(n1000));
  jnot g628(.din(n997), .dout(n1001));
  jor  g629(.dina(n678), .dinb(n909), .dout(n1002));
  jor  g630(.dina(n1002), .dinb(n1001), .dout(n1003));
  jand g631(.dina(n1003), .dinb(n1000), .dout(n1004));
  jxor g632(.dina(n716), .dinb(G1991), .dout(n1005));
  jor  g633(.dina(n1005), .dinb(n1001), .dout(n1006));
  jand g634(.dina(n1006), .dinb(n1004), .dout(n1007));
  jxor g635(.dina(n640), .dinb(n899), .dout(n1008));
  jxor g636(.dina(G290), .dinb(G1986), .dout(n1009));
  jand g637(.dina(n1009), .dinb(n1008), .dout(n1010));
  jor  g638(.dina(n1010), .dinb(n1001), .dout(n1011));
  jand g639(.dina(n1011), .dinb(n1007), .dout(n1012));
  jand g640(.dina(n1012), .dinb(n996), .dout(n1013));
  jnot g641(.din(G1986), .dout(n1014));
  jnot g642(.din(G290), .dout(n1015));
  jand g643(.dina(n1015), .dinb(n1014), .dout(n1016));
  jand g644(.dina(n1008), .dinb(n997), .dout(n1017));
  jand g645(.dina(n1017), .dinb(n1016), .dout(n1018));
  jand g646(.dina(n1018), .dinb(n1007), .dout(n1019));
  jnot g647(.din(n716), .dout(n1020));
  jand g648(.dina(n1020), .dinb(n610), .dout(n1021));
  jand g649(.dina(n1017), .dinb(n1021), .dout(n1022));
  jand g650(.dina(n1022), .dinb(n1004), .dout(n1023));
  jand g651(.dina(n640), .dinb(n899), .dout(n1024));
  jand g652(.dina(n1024), .dinb(n997), .dout(n1025));
  jand g653(.dina(n1025), .dinb(n1003), .dout(n1026));
  jor  g654(.dina(n1026), .dinb(n999), .dout(n1027));
  jor  g655(.dina(n1027), .dinb(n1023), .dout(n1028));
  jor  g656(.dina(n1028), .dinb(n1019), .dout(n1029));
  jor  g657(.dina(n1029), .dinb(n1013), .dout(G329));
  zero g658(.dout(G231));
  jor  g659(.dina(G229), .dinb(n503), .dout(n1032));
  jor  g660(.dina(n1032), .dinb(G227), .dout(n1033));
  jor  g661(.dina(n1033), .dinb(G401), .dout(n1034));
  jor  g662(.dina(n1034), .dinb(G397), .dout(n1035));
  jor  g663(.dina(n1035), .dinb(G395), .dout(G225));
  jnot g664(.din(G225), .dout(G308));
  buf  g665(.din(G452), .dout(G350));
  buf  g666(.din(G452), .dout(G335));
  buf  g667(.din(G452), .dout(G409));
  buf  g668(.din(G1083), .dout(G369));
  buf  g669(.din(G1083), .dout(G367));
  buf  g670(.din(G2066), .dout(G411));
  buf  g671(.din(G2066), .dout(G337));
  buf  g672(.din(G2066), .dout(G384));
  buf  g673(.din(G452), .dout(G391));
  jor  g674(.dina(n558), .dinb(n557), .dout(G321));
  jor  g675(.dina(n561), .dinb(n560), .dout(G280));
  jor  g676(.dina(n567), .dinb(n566), .dout(G323));
  jor  g677(.dina(n882), .dinb(n880), .dout(G331));
endmodule


